module Register #(parameter N = 32) (clk, In, Out);
    input clk;
    input [N-1:0] In, Out;
endmodule