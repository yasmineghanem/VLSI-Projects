module Radix4Booth ();
    
endmodule