module VerilogMultiplierTB ();
    
endmodule