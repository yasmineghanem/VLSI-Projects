module Radix4BoothTB ();
    
endmodule