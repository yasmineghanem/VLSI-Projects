module FLoatingPointMultiplierTB();
    
endmodule