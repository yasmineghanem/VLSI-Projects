module FLoatingPointMultiplier ();
    
endmodule