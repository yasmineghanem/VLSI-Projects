module BoothAlgorithm ();
    
endmodule