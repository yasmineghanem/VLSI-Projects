module MultiplierTreeTB ();
    
endmodule