module BoothAlgorithmTB ();
    
endmodule