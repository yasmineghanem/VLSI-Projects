module MultiplierTree ();
    
endmodule