module SequentialMultiplierTB();
    
endmodule