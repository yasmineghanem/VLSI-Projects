
// 	Wed Jan  4 11:26:31 2023
//	vlsi
//	localhost.localdomain

module datapath__0_253 (p_0, p_1);

output [63:0] p_1;
input [63:0] p_0;
wire slo__xsl_n176;
wire slo__sro_n91;
wire CLOCK_slo__sro_n317;
wire n_61;
wire n_0;
wire n_60;
wire n_59;
wire n_58;
wire n_57;
wire n_56;
wire n_55;
wire n_1;
wire n_54;
wire n_53;
wire n_52;
wire n_2;
wire n_51;
wire n_3;
wire n_50;
wire n_49;
wire n_47;
wire n_4;
wire n_48;
wire n_46;
wire n_5;
wire n_45;
wire n_44;
wire n_43;
wire n_42;
wire n_41;
wire n_40;
wire n_39;
wire n_38;
wire n_37;
wire n_36;
wire n_35;
wire n_34;
wire n_33;
wire n_32;
wire n_31;
wire n_30;
wire n_29;
wire n_28;
wire n_27;
wire n_26;
wire n_25;
wire n_24;
wire n_23;
wire n_22;
wire n_21;
wire n_20;
wire n_19;
wire n_18;
wire n_17;
wire n_16;
wire n_15;
wire n_14;
wire n_13;
wire n_12;
wire n_11;
wire n_6;
wire n_10;
wire n_9;
wire n_8;
wire n_7;
wire n_71;
wire n_70;
wire n_69;
wire n_68;
wire n_67;
wire n_66;
wire n_65;
wire n_64;
wire n_63;
wire n_62;
wire slo__n17;
wire slo__sro_n92;
wire CLOCK_slo__sro_n316;
wire slo__sro_n93;
wire slo__sro_n94;
wire CLOCK_slo__sro_n278;
wire CLOCK_slo__sro_n318;


INV_X4 i_134 (.ZN (n_71), .A (p_0[60]));
INV_X1 i_133 (.ZN (n_70), .A (p_0[55]));
INV_X1 i_132 (.ZN (n_69), .A (p_0[51]));
INV_X1 i_131 (.ZN (n_68), .A (p_0[45]));
INV_X1 i_130 (.ZN (n_67), .A (p_0[42]));
INV_X1 i_129 (.ZN (n_66), .A (p_0[36]));
INV_X1 i_128 (.ZN (n_65), .A (p_0[31]));
INV_X1 i_127 (.ZN (n_64), .A (p_0[27]));
INV_X1 i_126 (.ZN (n_63), .A (p_0[25]));
INV_X1 i_125 (.ZN (n_62), .A (p_0[6]));
OR3_X1 i_124 (.ZN (n_61), .A1 (p_0[2]), .A2 (p_0[1]), .A3 (p_0[0]));
OR2_X1 i_123 (.ZN (n_60), .A1 (n_61), .A2 (p_0[3]));
NOR2_X1 i_122 (.ZN (n_59), .A1 (n_60), .A2 (p_0[4]));
NOR3_X1 i_121 (.ZN (n_58), .A1 (n_60), .A2 (p_0[4]), .A3 (p_0[5]));
NAND2_X1 i_120 (.ZN (n_57), .A1 (n_58), .A2 (n_62));
OR2_X1 i_119 (.ZN (n_56), .A1 (n_57), .A2 (p_0[7]));
OR3_X1 i_118 (.ZN (n_55), .A1 (n_56), .A2 (p_0[8]), .A3 (p_0[9]));
OR2_X1 i_117 (.ZN (n_54), .A1 (n_55), .A2 (p_0[10]));
OR2_X1 i_116 (.ZN (n_53), .A1 (n_54), .A2 (p_0[11]));
OR3_X1 i_115 (.ZN (n_52), .A1 (n_53), .A2 (p_0[12]), .A3 (p_0[13]));
OR3_X2 i_114 (.ZN (n_51), .A1 (n_52), .A2 (p_0[14]), .A3 (p_0[15]));
OR2_X1 i_113 (.ZN (n_50), .A1 (n_51), .A2 (p_0[16]));
OR2_X1 i_112 (.ZN (n_49), .A1 (n_50), .A2 (p_0[17]));
NOR3_X2 i_111 (.ZN (n_48), .A1 (n_49), .A2 (p_0[18]), .A3 (p_0[19]));
INV_X2 i_110 (.ZN (n_47), .A (n_48));
OR3_X2 i_109 (.ZN (n_46), .A1 (n_47), .A2 (p_0[20]), .A3 (p_0[21]));
OR2_X1 i_108 (.ZN (n_45), .A1 (n_46), .A2 (p_0[22]));
NOR2_X1 i_107 (.ZN (n_44), .A1 (n_45), .A2 (p_0[23]));
NOR3_X1 i_106 (.ZN (n_43), .A1 (n_45), .A2 (p_0[23]), .A3 (p_0[24]));
NAND2_X1 i_105 (.ZN (n_42), .A1 (n_43), .A2 (n_63));
NOR2_X1 i_104 (.ZN (n_41), .A1 (n_42), .A2 (p_0[26]));
NAND2_X1 i_103 (.ZN (n_40), .A1 (n_41), .A2 (n_64));
NOR2_X1 i_102 (.ZN (n_39), .A1 (n_40), .A2 (p_0[28]));
NOR3_X1 i_101 (.ZN (n_38), .A1 (n_40), .A2 (p_0[28]), .A3 (p_0[29]));
NOR4_X2 i_100 (.ZN (n_37), .A1 (n_40), .A2 (p_0[28]), .A3 (p_0[29]), .A4 (p_0[30]));
NAND2_X1 i_99 (.ZN (n_36), .A1 (n_37), .A2 (n_65));
OR2_X1 i_98 (.ZN (n_35), .A1 (n_36), .A2 (p_0[32]));
NOR2_X1 i_97 (.ZN (n_34), .A1 (n_35), .A2 (p_0[33]));
NOR3_X1 i_96 (.ZN (n_33), .A1 (n_35), .A2 (p_0[33]), .A3 (p_0[34]));
NOR4_X4 i_95 (.ZN (n_32), .A1 (n_35), .A2 (p_0[33]), .A3 (p_0[34]), .A4 (p_0[35]));
NAND2_X1 i_94 (.ZN (n_31), .A1 (n_32), .A2 (n_66));
OR2_X1 i_93 (.ZN (n_30), .A1 (n_31), .A2 (p_0[37]));
OR2_X1 i_92 (.ZN (n_29), .A1 (n_30), .A2 (p_0[38]));
NOR2_X1 i_91 (.ZN (n_28), .A1 (n_29), .A2 (p_0[39]));
NOR3_X1 i_90 (.ZN (n_27), .A1 (n_29), .A2 (p_0[39]), .A3 (p_0[40]));
NOR4_X4 i_89 (.ZN (n_26), .A1 (p_0[41]), .A2 (p_0[39]), .A3 (p_0[40]), .A4 (n_29));
NAND2_X1 i_88 (.ZN (n_25), .A1 (n_26), .A2 (n_67));
NOR2_X2 i_87 (.ZN (n_24), .A1 (n_25), .A2 (p_0[43]));
NOR3_X1 i_86 (.ZN (n_23), .A1 (n_25), .A2 (p_0[43]), .A3 (p_0[44]));
NAND2_X1 i_85 (.ZN (n_22), .A1 (n_23), .A2 (n_68));
OR2_X1 i_84 (.ZN (n_21), .A1 (n_22), .A2 (p_0[46]));
OR2_X2 i_83 (.ZN (n_20), .A1 (n_21), .A2 (p_0[47]));
NOR2_X1 i_82 (.ZN (n_19), .A1 (n_20), .A2 (p_0[48]));
NOR3_X1 i_81 (.ZN (n_18), .A1 (n_20), .A2 (p_0[48]), .A3 (p_0[49]));
NOR4_X4 i_80 (.ZN (n_17), .A1 (n_20), .A2 (p_0[48]), .A3 (p_0[49]), .A4 (p_0[50]));
NAND2_X1 i_79 (.ZN (n_16), .A1 (n_17), .A2 (n_69));
NOR2_X1 i_78 (.ZN (n_15), .A1 (n_16), .A2 (p_0[52]));
NOR3_X1 i_77 (.ZN (n_14), .A1 (n_16), .A2 (p_0[52]), .A3 (p_0[53]));
NOR4_X4 i_76 (.ZN (n_13), .A1 (p_0[54]), .A2 (p_0[52]), .A3 (p_0[53]), .A4 (n_16));
NAND2_X1 i_75 (.ZN (n_12), .A1 (n_13), .A2 (n_70));
INV_X1 slo__xsl_c212 (.ZN (slo__xsl_n176), .A (slo__n17));
NOR2_X1 i_73 (.ZN (n_10), .A1 (slo__xsl_n176), .A2 (p_0[58]));
NOR3_X2 i_72 (.ZN (n_9), .A1 (p_0[59]), .A2 (p_0[58]), .A3 (slo__xsl_n176));
NAND2_X4 slo__sro_c124 (.ZN (slo__sro_n92), .A1 (slo__sro_n94), .A2 (slo__sro_n93));
NOR2_X4 i_70 (.ZN (n_7), .A1 (n_8), .A2 (p_0[61]));
INV_X4 slo__sro_c122 (.ZN (slo__sro_n94), .A (p_0[58]));
XNOR2_X2 i_68 (.ZN (p_1[62]), .A (p_0[62]), .B (n_7));
INV_X1 CLOCK_slo__sro_c360 (.ZN (CLOCK_slo__sro_n317), .A (n_12));
XNOR2_X1 i_66 (.ZN (p_1[60]), .A (p_0[60]), .B (n_9));
XNOR2_X1 i_65 (.ZN (p_1[59]), .A (p_0[59]), .B (n_10));
XOR2_X1 i_64 (.Z (p_1[58]), .A (p_0[58]), .B (slo__xsl_n176));
OAI21_X1 i_63 (.ZN (n_6), .A (p_0[57]), .B1 (n_12), .B2 (p_0[56]));
AND2_X1 i_62 (.ZN (p_1[57]), .A1 (slo__xsl_n176), .A2 (n_6));
XOR2_X1 i_61 (.Z (p_1[56]), .A (p_0[56]), .B (n_12));
XNOR2_X1 i_60 (.ZN (p_1[55]), .A (p_0[55]), .B (n_13));
XNOR2_X1 i_59 (.ZN (p_1[54]), .A (p_0[54]), .B (n_14));
XNOR2_X1 i_58 (.ZN (p_1[53]), .A (p_0[53]), .B (n_15));
XOR2_X1 i_57 (.Z (p_1[52]), .A (p_0[52]), .B (n_16));
XNOR2_X1 i_56 (.ZN (p_1[51]), .A (p_0[51]), .B (n_17));
XNOR2_X1 i_55 (.ZN (p_1[50]), .A (p_0[50]), .B (n_18));
XNOR2_X1 i_54 (.ZN (p_1[49]), .A (p_0[49]), .B (n_19));
XOR2_X1 i_53 (.Z (p_1[48]), .A (p_0[48]), .B (n_20));
XOR2_X1 i_52 (.Z (p_1[47]), .A (p_0[47]), .B (n_21));
XOR2_X1 i_51 (.Z (p_1[46]), .A (p_0[46]), .B (n_22));
XNOR2_X1 i_50 (.ZN (p_1[45]), .A (p_0[45]), .B (n_23));
XNOR2_X1 i_49 (.ZN (p_1[44]), .A (p_0[44]), .B (n_24));
XOR2_X1 i_48 (.Z (p_1[43]), .A (p_0[43]), .B (n_25));
XNOR2_X1 i_47 (.ZN (p_1[42]), .A (p_0[42]), .B (n_26));
XNOR2_X1 i_46 (.ZN (p_1[41]), .A (p_0[41]), .B (n_27));
XNOR2_X1 i_45 (.ZN (p_1[40]), .A (p_0[40]), .B (n_28));
XOR2_X1 i_44 (.Z (p_1[39]), .A (p_0[39]), .B (n_29));
XOR2_X1 i_43 (.Z (p_1[38]), .A (p_0[38]), .B (n_30));
XOR2_X1 i_42 (.Z (p_1[37]), .A (p_0[37]), .B (n_31));
XNOR2_X1 i_41 (.ZN (p_1[36]), .A (p_0[36]), .B (n_32));
XNOR2_X2 i_40 (.ZN (p_1[35]), .A (p_0[35]), .B (n_33));
XNOR2_X1 i_39 (.ZN (p_1[34]), .A (p_0[34]), .B (n_34));
XOR2_X1 i_38 (.Z (p_1[33]), .A (p_0[33]), .B (n_35));
XOR2_X1 i_37 (.Z (p_1[32]), .A (p_0[32]), .B (n_36));
XNOR2_X1 i_36 (.ZN (p_1[31]), .A (p_0[31]), .B (n_37));
XNOR2_X1 i_35 (.ZN (p_1[30]), .A (p_0[30]), .B (n_38));
XNOR2_X1 i_34 (.ZN (p_1[29]), .A (p_0[29]), .B (n_39));
XOR2_X1 i_33 (.Z (p_1[28]), .A (p_0[28]), .B (n_40));
XNOR2_X1 i_32 (.ZN (p_1[27]), .A (p_0[27]), .B (n_41));
XOR2_X1 i_31 (.Z (p_1[26]), .A (p_0[26]), .B (n_42));
XNOR2_X1 i_30 (.ZN (p_1[25]), .A (p_0[25]), .B (n_43));
XNOR2_X1 i_29 (.ZN (p_1[24]), .A (p_0[24]), .B (n_44));
XOR2_X1 i_28 (.Z (p_1[23]), .A (p_0[23]), .B (n_45));
XOR2_X1 i_27 (.Z (p_1[22]), .A (p_0[22]), .B (n_46));
OAI21_X1 i_26 (.ZN (n_5), .A (p_0[21]), .B1 (n_47), .B2 (p_0[20]));
AND2_X1 i_25 (.ZN (p_1[21]), .A1 (n_46), .A2 (n_5));
XNOR2_X1 i_24 (.ZN (p_1[20]), .A (p_0[20]), .B (n_48));
OAI21_X1 i_23 (.ZN (n_4), .A (p_0[19]), .B1 (n_49), .B2 (p_0[18]));
AND2_X1 i_22 (.ZN (p_1[19]), .A1 (n_47), .A2 (n_4));
XOR2_X1 i_21 (.Z (p_1[18]), .A (p_0[18]), .B (n_49));
XOR2_X1 i_20 (.Z (p_1[17]), .A (p_0[17]), .B (n_50));
XOR2_X1 i_19 (.Z (p_1[16]), .A (p_0[16]), .B (n_51));
OAI21_X1 i_18 (.ZN (n_3), .A (p_0[15]), .B1 (n_52), .B2 (p_0[14]));
AND2_X1 i_17 (.ZN (p_1[15]), .A1 (n_51), .A2 (n_3));
XOR2_X1 i_16 (.Z (p_1[14]), .A (p_0[14]), .B (n_52));
OAI21_X1 i_15 (.ZN (n_2), .A (p_0[13]), .B1 (n_53), .B2 (p_0[12]));
AND2_X1 i_14 (.ZN (p_1[13]), .A1 (n_52), .A2 (n_2));
XOR2_X1 i_13 (.Z (p_1[12]), .A (p_0[12]), .B (n_53));
XOR2_X1 i_12 (.Z (p_1[11]), .A (p_0[11]), .B (n_54));
XOR2_X1 i_11 (.Z (p_1[10]), .A (p_0[10]), .B (n_55));
OAI21_X1 i_10 (.ZN (n_1), .A (p_0[9]), .B1 (n_56), .B2 (p_0[8]));
AND2_X1 i_9 (.ZN (p_1[9]), .A1 (n_55), .A2 (n_1));
XOR2_X1 i_8 (.Z (p_1[8]), .A (p_0[8]), .B (n_56));
XOR2_X1 i_7 (.Z (p_1[7]), .A (p_0[7]), .B (n_57));
XNOR2_X1 i_6 (.ZN (p_1[6]), .A (p_0[6]), .B (n_58));
XNOR2_X1 i_5 (.ZN (p_1[5]), .A (p_0[5]), .B (n_59));
XOR2_X1 i_4 (.Z (p_1[4]), .A (p_0[4]), .B (n_60));
XOR2_X1 i_3 (.Z (p_1[3]), .A (p_0[3]), .B (n_61));
OAI21_X1 i_2 (.ZN (n_0), .A (p_0[2]), .B1 (p_0[1]), .B2 (p_0[0]));
AND2_X1 i_1 (.ZN (p_1[2]), .A1 (n_61), .A2 (n_0));
XOR2_X1 i_0 (.Z (p_1[1]), .A (p_0[1]), .B (p_0[0]));
INV_X1 slo__c40 (.ZN (n_11), .A (slo__n17));
INV_X4 CLOCK_slo__sro_c359 (.ZN (CLOCK_slo__sro_n318), .A (p_0[56]));
NOR2_X1 slo__mro_c52 (.ZN (p_1[63]), .A1 (p_0[62]), .A2 (n_7));
INV_X2 slo__sro_c123 (.ZN (slo__sro_n93), .A (n_11));
INV_X2 CLOCK_slo__sro_c326 (.ZN (CLOCK_slo__sro_n278), .A (n_8));
NAND2_X4 slo__sro_c89 (.ZN (n_8), .A1 (n_71), .A2 (slo__sro_n91));
NOR2_X4 slo__sro_c125 (.ZN (slo__sro_n91), .A1 (p_0[59]), .A2 (slo__sro_n92));
XNOR2_X2 CLOCK_slo__sro_c327 (.ZN (p_1[61]), .A (p_0[61]), .B (CLOCK_slo__sro_n278));
NAND2_X2 CLOCK_slo__sro_c361 (.ZN (CLOCK_slo__sro_n316), .A1 (CLOCK_slo__sro_n317), .A2 (CLOCK_slo__sro_n318));
NOR2_X4 CLOCK_slo__sro_c362 (.ZN (slo__n17), .A1 (CLOCK_slo__sro_n316), .A2 (p_0[57]));

endmodule //datapath__0_253

module datapath__0_247 (p_1_25_PP_0, p_1_25_PP_1, p_0, p_1, p_2);

output [31:0] p_2;
input [31:0] p_0;
input [31:0] p_1;
input p_1_25_PP_0;
input p_1_25_PP_1;
wire n_1;
wire n_2;
wire n_3;
wire n_4;
wire n_5;
wire n_6;
wire n_7;
wire n_8;
wire n_10;
wire n_11;
wire n_12;
wire n_13;
wire n_14;
wire n_15;
wire n_16;
wire n_17;
wire slo__sro_n682;
wire n_19;
wire slo__sro_n436;
wire n_21;
wire slo__sro_n258;
wire n_24;
wire n_25;
wire n_28;
wire n_32;
wire n_0;
wire n_34;
wire n_33;
wire sgo__sro_n61;
wire sgo__sro_n62;
wire sgo__sro_n63;
wire sgo__sro_n64;
wire sgo__sro_n65;
wire sgo__sro_n66;
wire sgo__sro_n67;
wire slo__sro_n97;
wire slo__sro_n98;
wire slo__sro_n99;
wire slo__sro_n100;
wire slo__sro_n116;
wire slo__sro_n117;
wire slo__sro_n119;
wire slo__sro_n120;
wire slo__sro_n121;
wire slo__sro_n122;
wire slo__sro_n137;
wire slo__sro_n138;
wire slo__sro_n139;
wire slo__sro_n140;
wire slo__sro_n141;
wire slo__sro_n156;
wire slo__sro_n157;
wire slo__sro_n158;
wire slo__sro_n159;
wire slo__sro_n160;
wire slo__sro_n162;
wire slo__sro_n189;
wire slo__sro_n190;
wire slo__sro_n191;
wire slo__sro_n192;
wire slo__n415;
wire slo__sro_n255;
wire slo__sro_n256;
wire slo__sro_n257;
wire slo__sro_n217;
wire slo__sro_n218;
wire slo__sro_n219;
wire slo__sro_n220;
wire slo__sro_n221;
wire slo__sro_n275;
wire slo__sro_n276;
wire slo__sro_n277;
wire slo__sro_n278;
wire slo__sro_n434;
wire slo__sro_n435;
wire slo__sro_n365;
wire slo__sro_n366;
wire slo__sro_n367;
wire slo__sro_n368;
wire slo__sro_n369;
wire slo__sro_n437;
wire slo__sro_n438;
wire slo__sro_n439;
wire slo__sro_n681;
wire slo__sro_n604;
wire slo__sro_n605;
wire slo__sro_n606;
wire slo__sro_n607;
wire slo__sro_n608;
wire slo__sro_n609;
wire slo__sro_n610;
wire slo__sro_n683;
wire slo__sro_n684;
wire slo__sro_n863;
wire slo__sro_n864;
wire slo__sro_n796;
wire slo__sro_n860;
wire slo__sro_n861;
wire slo__sro_n862;
wire CLOCK_slo__sro_n1598;
wire CLOCK_slo__sro_n1599;
wire CLOCK_slo__sro_n1600;
wire CLOCK_slo__sro_n1601;
wire CLOCK_slo__sro_n1648;
wire CLOCK_slo__sro_n1649;
wire CLOCK_slo__sro_n1650;
wire CLOCK_slo__sro_n1651;
wire CLOCK_slo__sro_n1699;
wire CLOCK_slo__sro_n1700;
wire CLOCK_slo__sro_n1701;
wire CLOCK_slo__sro_n1702;
wire CLOCK_slo__sro_n1712;
wire CLOCK_slo__sro_n1713;
wire CLOCK_slo__sro_n1714;
wire CLOCK_slo__sro_n1715;
wire CLOCK_slo__xsl_n1987;
wire CLOCK_slo__sro_n1882;


INV_X1 i_36 (.ZN (n_34), .A (p_0[30]));
INV_X1 i_35 (.ZN (n_33), .A (p_1[30]));
INV_X1 i_34 (.ZN (n_32), .A (slo__sro_n98));
XNOR2_X1 slo__sro_c600 (.ZN (p_2[28]), .A (n_28), .B (slo__sro_n116));
OAI22_X1 i_31 (.ZN (n_0), .A1 (n_34), .A2 (p_1[30]), .B1 (p_0[30]), .B2 (n_33));
XNOR2_X1 i_0 (.ZN (p_2[30]), .A (n_32), .B (n_0));
INV_X1 slo__sro_c52 (.ZN (slo__sro_n122), .A (p_0[28]));
INV_X2 slo__sro_c70 (.ZN (slo__sro_n141), .A (slo__sro_n157));
FA_X1 i_28 (.CO (n_28), .S (p_2[27]), .A (p_0[27]), .B (p_1[27]), .CI (slo__sro_n138));
INV_X1 slo__sro_c86 (.ZN (slo__sro_n162), .A (p_0[25]));
INV_X1 slo__sro_c117 (.ZN (slo__sro_n192), .A (n_4));
FA_X1 i_25 (.CO (n_25), .S (p_2[24]), .A (p_0[24]), .B (p_1[24]), .CI (n_24));
FA_X1 i_24 (.CO (n_24), .S (p_2[23]), .A (p_0[23]), .B (p_1[23]), .CI (CLOCK_slo__sro_n1713));
XNOR2_X1 slo__sro_c177 (.ZN (slo__sro_n255), .A (p_1[3]), .B (p_0[3]));
NAND2_X1 slo__sro_c323 (.ZN (slo__sro_n436), .A1 (slo__sro_n438), .A2 (slo__sro_n439));
NAND2_X1 slo__sro_c501 (.ZN (slo__sro_n683), .A1 (p_1[9]), .A2 (p_0[9]));
NOR2_X4 slo__sro_c502 (.ZN (slo__sro_n682), .A1 (p_1[9]), .A2 (p_0[9]));
INV_X2 CLOCK_slo__sro_c1365 (.ZN (CLOCK_slo__sro_n1651), .A (n_15));
FA_X1 i_15 (.CO (n_15), .S (p_2[14]), .A (p_0[14]), .B (p_1[14]), .CI (n_14));
FA_X1 i_14 (.CO (n_14), .S (p_2[13]), .A (p_0[13]), .B (p_1[13]), .CI (n_13));
FA_X1 i_13 (.CO (n_13), .S (p_2[12]), .A (p_0[12]), .B (p_1[12]), .CI (n_12));
FA_X1 i_12 (.CO (n_12), .S (p_2[11]), .A (p_0[11]), .B (p_1[11]), .CI (n_11));
FA_X1 i_11 (.CO (n_11), .S (p_2[10]), .A (p_0[10]), .B (p_1[10]), .CI (n_10));
INV_X1 slo__sro_c594 (.ZN (slo__sro_n796), .A (p_0[31]));
NAND2_X1 CLOCK_slo__sro_c1432 (.ZN (CLOCK_slo__sro_n1715), .A1 (p_0[22]), .A2 (slo__sro_n218));
FA_X1 i_7 (.CO (n_7), .S (p_2[6]), .A (p_0[6]), .B (p_1[6]), .CI (n_6));
FA_X1 i_6 (.CO (n_6), .S (p_2[5]), .A (p_0[5]), .B (p_1[5]), .CI (n_5));
INV_X1 slo__sro_c320 (.ZN (slo__sro_n439), .A (p_0[18]));
INV_X2 slo__sro_c194 (.ZN (slo__sro_n278), .A (slo__n415));
FA_X1 i_3 (.CO (n_3), .S (p_2[2]), .A (p_0[2]), .B (p_1[2]), .CI (n_2));
FA_X1 i_2 (.CO (n_2), .S (p_2[1]), .A (p_0[1]), .B (p_1[1]), .CI (n_1));
HA_X1 i_1 (.CO (n_1), .S (p_2[0]), .A (p_0[0]), .B (p_1[0]));
INV_X1 sgo__sro_c1 (.ZN (sgo__sro_n67), .A (n_34));
INV_X1 sgo__sro_c2 (.ZN (sgo__sro_n66), .A (p_1[30]));
INV_X1 sgo__sro_c3 (.ZN (sgo__sro_n65), .A (p_0[30]));
INV_X1 sgo__sro_c4 (.ZN (sgo__sro_n64), .A (n_33));
NAND2_X1 sgo__sro_c5 (.ZN (sgo__sro_n63), .A1 (sgo__sro_n64), .A2 (sgo__sro_n65));
NAND2_X1 sgo__sro_c6 (.ZN (sgo__sro_n62), .A1 (sgo__sro_n66), .A2 (sgo__sro_n67));
OAI22_X1 sgo__sro_c7 (.ZN (sgo__sro_n61), .A1 (slo__sro_n98), .A2 (sgo__sro_n63), .B1 (n_32), .B2 (sgo__sro_n62));
NAND2_X1 slo__sro_c37 (.ZN (slo__sro_n100), .A1 (p_1[29]), .A2 (p_0[29]));
NOR2_X2 slo__sro_c38 (.ZN (slo__sro_n99), .A1 (p_1[29]), .A2 (p_0[29]));
OAI21_X2 slo__sro_c39 (.ZN (slo__sro_n98), .A (slo__sro_n100), .B1 (slo__sro_n117), .B2 (slo__sro_n99));
XNOR2_X1 slo__sro_c40 (.ZN (slo__sro_n97), .A (p_1[29]), .B (p_0[29]));
XNOR2_X2 slo__sro_c41 (.ZN (p_2[29]), .A (CLOCK_slo__xsl_n1987), .B (slo__sro_n97));
INV_X1 slo__sro_c53 (.ZN (slo__sro_n121), .A (p_1[28]));
NAND2_X1 slo__sro_c54 (.ZN (slo__sro_n120), .A1 (p_1[28]), .A2 (p_0[28]));
NAND2_X1 slo__sro_c55 (.ZN (slo__sro_n119), .A1 (slo__sro_n121), .A2 (slo__sro_n122));
INV_X1 CLOCK_slo__xsl_c1717 (.ZN (CLOCK_slo__xsl_n1987), .A (slo__sro_n117));
XNOR2_X1 slo__sro_c58 (.ZN (slo__sro_n116), .A (p_1[28]), .B (p_0[28]));
INV_X1 slo__sro_c632 (.ZN (slo__sro_n864), .A (n_8));
NAND2_X1 slo__sro_c71 (.ZN (slo__sro_n140), .A1 (p_1[26]), .A2 (p_0[26]));
NOR2_X2 slo__sro_c72 (.ZN (slo__sro_n139), .A1 (p_1[26]), .A2 (p_0[26]));
OAI21_X2 slo__sro_c73 (.ZN (slo__sro_n138), .A (slo__sro_n140), .B1 (slo__sro_n141), .B2 (slo__sro_n139));
XNOR2_X1 slo__sro_c74 (.ZN (slo__sro_n137), .A (p_1[26]), .B (p_0[26]));
XNOR2_X1 slo__sro_c75 (.ZN (p_2[26]), .A (slo__sro_n137), .B (slo__sro_n157));
INV_X1 slo__sro_c500 (.ZN (slo__sro_n684), .A (slo__sro_n861));
NAND2_X1 slo__sro_c88 (.ZN (slo__sro_n160), .A1 (p_1_25_PP_0), .A2 (p_0[25]));
NAND2_X1 slo__sro_c89 (.ZN (slo__sro_n159), .A1 (p_1_25_PP_1), .A2 (slo__sro_n162));
NAND2_X2 slo__sro_c90 (.ZN (slo__sro_n158), .A1 (n_25), .A2 (slo__sro_n159));
NAND2_X2 slo__sro_c91 (.ZN (slo__sro_n157), .A1 (slo__sro_n158), .A2 (slo__sro_n160));
XNOR2_X1 slo__sro_c92 (.ZN (slo__sro_n156), .A (p_1[25]), .B (p_0[25]));
XNOR2_X1 slo__sro_c93 (.ZN (p_2[25]), .A (n_25), .B (slo__sro_n156));
NAND2_X1 slo__sro_c118 (.ZN (slo__sro_n191), .A1 (p_1[4]), .A2 (p_0[4]));
NOR2_X1 slo__sro_c119 (.ZN (slo__sro_n190), .A1 (p_1[4]), .A2 (p_0[4]));
OAI21_X1 slo__sro_c120 (.ZN (n_5), .A (slo__sro_n191), .B1 (slo__sro_n192), .B2 (slo__sro_n190));
XNOR2_X1 slo__sro_c121 (.ZN (slo__sro_n189), .A (p_1[4]), .B (p_0[4]));
XNOR2_X1 slo__sro_c122 (.ZN (p_2[4]), .A (slo__sro_n189), .B (n_4));
OAI21_X2 slo__c303 (.ZN (slo__n415), .A (slo__sro_n368), .B1 (slo__sro_n369), .B2 (slo__sro_n367));
INV_X1 slo__sro_c173 (.ZN (slo__sro_n258), .A (n_3));
NAND2_X1 slo__sro_c174 (.ZN (slo__sro_n257), .A1 (p_1[3]), .A2 (p_0[3]));
NOR2_X1 slo__sro_c175 (.ZN (slo__sro_n256), .A1 (p_1[3]), .A2 (p_0[3]));
OAI21_X1 slo__sro_c176 (.ZN (n_4), .A (slo__sro_n257), .B1 (slo__sro_n258), .B2 (slo__sro_n256));
INV_X2 slo__sro_c144 (.ZN (slo__sro_n221), .A (n_21));
NAND2_X1 slo__sro_c145 (.ZN (slo__sro_n220), .A1 (p_1[21]), .A2 (p_0[21]));
NOR2_X2 slo__sro_c146 (.ZN (slo__sro_n219), .A1 (p_1[21]), .A2 (p_0[21]));
OAI21_X2 slo__sro_c147 (.ZN (slo__sro_n218), .A (slo__sro_n220), .B1 (slo__sro_n221), .B2 (slo__sro_n219));
XNOR2_X1 slo__sro_c148 (.ZN (slo__sro_n217), .A (p_1[21]), .B (p_0[21]));
XNOR2_X1 slo__sro_c149 (.ZN (p_2[21]), .A (n_21), .B (slo__sro_n217));
XNOR2_X1 slo__sro_c178 (.ZN (p_2[3]), .A (slo__sro_n255), .B (n_3));
NAND2_X1 slo__sro_c195 (.ZN (slo__sro_n277), .A1 (p_1[20]), .A2 (p_0[20]));
NOR2_X4 slo__sro_c196 (.ZN (slo__sro_n276), .A1 (p_1[20]), .A2 (p_0[20]));
OAI21_X2 slo__sro_c197 (.ZN (n_21), .A (slo__sro_n277), .B1 (slo__sro_n278), .B2 (slo__sro_n276));
XNOR2_X1 slo__sro_c198 (.ZN (slo__sro_n275), .A (p_1[20]), .B (p_0[20]));
XNOR2_X1 slo__sro_c199 (.ZN (p_2[20]), .A (slo__sro_n366), .B (slo__sro_n275));
INV_X1 slo__sro_c321 (.ZN (slo__sro_n438), .A (p_1[18]));
NAND2_X1 slo__sro_c322 (.ZN (slo__sro_n437), .A1 (p_1[18]), .A2 (p_0[18]));
INV_X2 slo__sro_c272 (.ZN (slo__sro_n369), .A (n_19));
NAND2_X1 slo__sro_c273 (.ZN (slo__sro_n368), .A1 (p_1[19]), .A2 (p_0[19]));
NOR2_X1 slo__sro_c274 (.ZN (slo__sro_n367), .A1 (p_1[19]), .A2 (p_0[19]));
OAI21_X1 slo__sro_c275 (.ZN (slo__sro_n366), .A (slo__sro_n368), .B1 (slo__sro_n369), .B2 (slo__sro_n367));
XNOR2_X1 slo__sro_c276 (.ZN (slo__sro_n365), .A (p_1[19]), .B (p_0[19]));
XNOR2_X1 slo__sro_c277 (.ZN (p_2[19]), .A (n_19), .B (slo__sro_n365));
NAND2_X2 slo__sro_c324 (.ZN (slo__sro_n435), .A1 (slo__sro_n605), .A2 (slo__sro_n436));
NAND2_X2 slo__sro_c325 (.ZN (n_19), .A1 (slo__sro_n435), .A2 (slo__sro_n437));
XNOR2_X1 slo__sro_c326 (.ZN (slo__sro_n434), .A (p_1[18]), .B (p_0[18]));
XNOR2_X1 slo__sro_c327 (.ZN (p_2[18]), .A (slo__sro_n605), .B (slo__sro_n434));
INV_X1 slo__sro_c437 (.ZN (slo__sro_n610), .A (p_0[17]));
INV_X1 slo__sro_c438 (.ZN (slo__sro_n609), .A (p_1[17]));
NAND2_X1 slo__sro_c439 (.ZN (slo__sro_n608), .A1 (p_1[17]), .A2 (p_0[17]));
NAND2_X1 slo__sro_c440 (.ZN (slo__sro_n607), .A1 (slo__sro_n610), .A2 (slo__sro_n609));
NAND2_X2 slo__sro_c441 (.ZN (slo__sro_n606), .A1 (n_17), .A2 (slo__sro_n607));
NAND2_X2 slo__sro_c442 (.ZN (slo__sro_n605), .A1 (slo__sro_n606), .A2 (slo__sro_n608));
XNOR2_X1 slo__sro_c443 (.ZN (slo__sro_n604), .A (p_1[17]), .B (p_0[17]));
XNOR2_X1 slo__sro_c444 (.ZN (p_2[17]), .A (n_17), .B (slo__sro_n604));
OAI21_X1 slo__sro_c503 (.ZN (n_10), .A (slo__sro_n683), .B1 (slo__sro_n684), .B2 (slo__sro_n682));
XNOR2_X1 slo__sro_c504 (.ZN (slo__sro_n681), .A (p_1[9]), .B (p_0[9]));
XNOR2_X1 slo__sro_c505 (.ZN (p_2[9]), .A (slo__sro_n681), .B (slo__sro_n861));
XNOR2_X1 slo__sro_c595 (.ZN (p_2[31]), .A (sgo__sro_n61), .B (slo__sro_n796));
INV_X2 CLOCK_slo__sro_c1312 (.ZN (CLOCK_slo__sro_n1601), .A (n_16));
NAND2_X1 CLOCK_slo__sro_c1313 (.ZN (CLOCK_slo__sro_n1600), .A1 (p_1[16]), .A2 (p_0[16]));
NAND2_X1 slo__sro_c633 (.ZN (slo__sro_n863), .A1 (p_1[8]), .A2 (p_0[8]));
NOR2_X1 slo__sro_c634 (.ZN (slo__sro_n862), .A1 (p_1[8]), .A2 (p_0[8]));
OAI21_X2 slo__sro_c635 (.ZN (slo__sro_n861), .A (slo__sro_n863), .B1 (slo__sro_n864), .B2 (slo__sro_n862));
XNOR2_X1 slo__sro_c636 (.ZN (slo__sro_n860), .A (p_1[8]), .B (p_0[8]));
XNOR2_X1 slo__sro_c637 (.ZN (p_2[8]), .A (slo__sro_n860), .B (n_8));
NOR2_X1 CLOCK_slo__sro_c1314 (.ZN (CLOCK_slo__sro_n1599), .A1 (p_1[16]), .A2 (p_0[16]));
OAI21_X4 CLOCK_slo__sro_c1315 (.ZN (n_17), .A (CLOCK_slo__sro_n1600), .B1 (CLOCK_slo__sro_n1601), .B2 (CLOCK_slo__sro_n1599));
XNOR2_X1 CLOCK_slo__sro_c1316 (.ZN (CLOCK_slo__sro_n1598), .A (p_1[16]), .B (p_0[16]));
XNOR2_X1 CLOCK_slo__sro_c1317 (.ZN (p_2[16]), .A (n_16), .B (CLOCK_slo__sro_n1598));
NAND2_X1 CLOCK_slo__sro_c1366 (.ZN (CLOCK_slo__sro_n1650), .A1 (p_1[15]), .A2 (p_0[15]));
NOR2_X2 CLOCK_slo__sro_c1367 (.ZN (CLOCK_slo__sro_n1649), .A1 (p_1[15]), .A2 (p_0[15]));
OAI21_X2 CLOCK_slo__sro_c1368 (.ZN (n_16), .A (CLOCK_slo__sro_n1650), .B1 (CLOCK_slo__sro_n1651), .B2 (CLOCK_slo__sro_n1649));
XNOR2_X1 CLOCK_slo__sro_c1369 (.ZN (CLOCK_slo__sro_n1648), .A (p_1[15]), .B (p_0[15]));
XNOR2_X1 CLOCK_slo__sro_c1370 (.ZN (p_2[15]), .A (n_15), .B (CLOCK_slo__sro_n1648));
INV_X2 CLOCK_slo__sro_c1418 (.ZN (CLOCK_slo__sro_n1702), .A (n_7));
NAND2_X1 CLOCK_slo__sro_c1419 (.ZN (CLOCK_slo__sro_n1701), .A1 (p_1[7]), .A2 (p_0[7]));
NOR2_X2 CLOCK_slo__sro_c1420 (.ZN (CLOCK_slo__sro_n1700), .A1 (p_1[7]), .A2 (p_0[7]));
OAI21_X4 CLOCK_slo__sro_c1421 (.ZN (n_8), .A (CLOCK_slo__sro_n1701), .B1 (CLOCK_slo__sro_n1702), .B2 (CLOCK_slo__sro_n1700));
XNOR2_X1 CLOCK_slo__sro_c1422 (.ZN (CLOCK_slo__sro_n1699), .A (p_1[7]), .B (p_0[7]));
XNOR2_X1 CLOCK_slo__sro_c1423 (.ZN (p_2[7]), .A (CLOCK_slo__sro_n1699), .B (n_7));
AOI22_X2 CLOCK_slo__sro_c1433 (.ZN (CLOCK_slo__sro_n1714), .A1 (slo__sro_n218), .A2 (p_1[22])
    , .B1 (p_1[22]), .B2 (p_0[22]));
NAND2_X2 CLOCK_slo__sro_c1434 (.ZN (CLOCK_slo__sro_n1713), .A1 (CLOCK_slo__sro_n1714), .A2 (CLOCK_slo__sro_n1715));
XNOR2_X1 CLOCK_slo__sro_c1435 (.ZN (CLOCK_slo__sro_n1712), .A (p_1[22]), .B (p_0[22]));
XNOR2_X1 CLOCK_slo__sro_c1436 (.ZN (p_2[22]), .A (CLOCK_slo__sro_n1712), .B (slo__sro_n218));
NAND2_X2 CLOCK_slo__sro_c1605 (.ZN (CLOCK_slo__sro_n1882), .A1 (n_28), .A2 (slo__sro_n119));
AND2_X4 CLOCK_slo__xsl_c1720 (.ZN (slo__sro_n117), .A1 (CLOCK_slo__sro_n1882), .A2 (slo__sro_n120));

endmodule //datapath__0_247

module datapath__0_246 (drc_ipoPP_0, Multiplier, p_0, p_1);

output [31:0] p_1;
input [31:0] Multiplier;
input [31:0] p_0;
input drc_ipoPP_0;
wire slo__n353;
wire n_1;
wire n_2;
wire n_3;
wire n_4;
wire CLOCK_slo__xsl_n1571;
wire n_6;
wire n_7;
wire n_8;
wire n_9;
wire n_10;
wire n_11;
wire n_12;
wire n_14;
wire slo__sro_n180;
wire n_16;
wire n_17;
wire n_18;
wire n_19;
wire n_21;
wire n_22;
wire n_23;
wire n_24;
wire slo__xsl_n847;
wire CLOCK_slo__sro_n1252;
wire n_27;
wire n_28;
wire n_0;
wire n_34;
wire n_33;
wire sgo__sro_n57;
wire sgo__sro_n58;
wire CLOCK_slo__sro_n1251;
wire sgo__sro_n60;
wire slo__xsl_n846;
wire slo__sro_n85;
wire slo__sro_n86;
wire slo__sro_n87;
wire slo__sro_n88;
wire slo__sro_n89;
wire slo__sro_n106;
wire slo__sro_n107;
wire slo__sro_n108;
wire slo__sro_n109;
wire slo__sro_n159;
wire slo__sro_n160;
wire slo__sro_n161;
wire slo__sro_n162;
wire slo__sro_n163;
wire slo__sro_n134;
wire slo__sro_n135;
wire slo__sro_n136;
wire slo__sro_n137;
wire slo__sro_n138;
wire slo__sro_n181;
wire slo__sro_n182;
wire slo__sro_n183;
wire slo__sro_n199;
wire slo__sro_n200;
wire slo__sro_n201;
wire slo__sro_n202;
wire slo__sro_n203;
wire slo__sro_n219;
wire slo__sro_n220;
wire slo__sro_n221;
wire slo__sro_n222;
wire slo__sro_n232;
wire slo__sro_n233;
wire slo__sro_n234;
wire slo__sro_n235;
wire slo__sro_n236;
wire slo__sro_n591;
wire slo__n313;
wire slo__n401;
wire slo__sro_n328;
wire slo__sro_n453;
wire slo__sro_n454;
wire slo__sro_n455;
wire slo__sro_n456;
wire slo__n531;
wire slo__sro_n592;
wire slo__sro_n593;
wire slo__sro_n594;
wire slo__sro_n595;
wire slo__sro_n596;
wire slo__sro_n768;
wire slo__sro_n769;
wire opt_ipo_n619;
wire slo__sro_n734;
wire slo__sro_n735;
wire slo__sro_n736;
wire slo__sro_n737;
wire slo__sro_n770;
wire slo__sro_n771;
wire slo__sro_n772;
wire slo__sro_n785;
wire slo__sro_n786;
wire slo__sro_n787;
wire slo__sro_n788;
wire slo__sro_n789;
wire CLOCK_slo__sro_n1250;
wire slo__mro_n810;
wire CLOCK_slo__sro_n1249;
wire CLOCK_slo__sro_n1315;
wire CLOCK_slo__sro_n1316;
wire CLOCK_slo__sro_n1317;
wire CLOCK_slo__sro_n1318;
wire CLOCK_slo__sro_n1414;
wire CLOCK_slo__sro_n1415;
wire CLOCK_slo__sro_n1416;
wire CLOCK_slo__sro_n1417;
wire CLOCK_slo__sro_n1446;
wire CLOCK_slo__xsl_n1572;
wire CLOCK_slo__sro_n1622;
wire CLOCK_slo__xsl_n1478;
wire CLOCK_slo__xsl_n1479;
wire CLOCK_slo__sro_n1623;
wire CLOCK_slo__sro_n1624;
wire CLOCK_slo__sro_n1625;


INV_X1 i_36 (.ZN (n_34), .A (Multiplier[30]));
INV_X2 i_35 (.ZN (n_33), .A (p_0[30]));
INV_X2 slo__sro_c599 (.ZN (slo__sro_n737), .A (n_17));
INV_X2 slo__sro_c29 (.ZN (slo__sro_n89), .A (slo__sro_n160));
OAI21_X1 slo__c312 (.ZN (slo__n401), .A (slo__sro_n221), .B1 (slo__sro_n222), .B2 (slo__sro_n220));
OAI22_X1 i_31 (.ZN (n_0), .A1 (n_34), .A2 (p_0[30]), .B1 (n_33), .B2 (Multiplier[30]));
XNOR2_X1 i_0 (.ZN (p_1[30]), .A (n_0), .B (opt_ipo_n619));
INV_X1 slo__sro_c50 (.ZN (slo__sro_n109), .A (n_4));
INV_X1 slo__sro_c120 (.ZN (slo__sro_n183), .A (n_27));
INV_X1 slo__sro_c143 (.ZN (slo__sro_n203), .A (slo__n401));
INV_X1 slo__xsl_c686 (.ZN (slo__xsl_n846), .A (slo__xsl_n847));
OAI21_X1 slo__c402 (.ZN (slo__n531), .A (slo__sro_n455), .B1 (slo__sro_n456), .B2 (slo__sro_n454));
INV_X2 CLOCK_slo__sro_c1047 (.ZN (CLOCK_slo__sro_n1318), .A (n_11));
FA_X1 i_22 (.CO (n_22), .S (p_1[21]), .A (Multiplier[21]), .B (p_0[21]), .CI (n_21));
FA_X1 i_21 (.CO (n_21), .S (p_1[20]), .A (Multiplier[20]), .B (p_0[20]), .CI (slo__sro_n200));
INV_X2 slo__sro_c160 (.ZN (slo__sro_n222), .A (n_18));
INV_X1 slo__sro_c174 (.ZN (slo__sro_n236), .A (slo__n531));
INV_X2 slo__sro_c622 (.ZN (slo__sro_n772), .A (n_12));
FA_X1 i_17 (.CO (n_17), .S (p_1[16]), .A (Multiplier[16]), .B (p_0[16]), .CI (n_16));
OAI21_X2 CLOCK_slo__sro_c1188 (.ZN (CLOCK_slo__sro_n1446), .A (slo__sro_n108), .B1 (slo__sro_n109), .B2 (slo__sro_n107));
NAND2_X1 slo__sro_c121 (.ZN (slo__sro_n182), .A1 (p_0[27]), .A2 (Multiplier[27]));
NOR2_X1 slo__sro_c624 (.ZN (slo__sro_n770), .A1 (p_0[12]), .A2 (Multiplier[12]));
INV_X1 slo__sro_c636 (.ZN (slo__sro_n789), .A (slo__sro_n233));
INV_X2 CLOCK_slo__sro_c1157 (.ZN (CLOCK_slo__sro_n1417), .A (slo__sro_n135));
FA_X1 i_11 (.CO (n_11), .S (p_1[10]), .A (Multiplier[10]), .B (p_0[10]), .CI (n_10));
FA_X1 i_10 (.CO (n_10), .S (p_1[9]), .A (Multiplier[9]), .B (p_0[9]), .CI (n_9));
FA_X1 i_9 (.CO (n_9), .S (p_1[8]), .A (Multiplier[8]), .B (p_0[8]), .CI (n_8));
FA_X1 i_8 (.CO (n_8), .S (p_1[7]), .A (Multiplier[7]), .B (p_0[7]), .CI (n_7));
FA_X1 i_7 (.CO (n_7), .S (p_1[6]), .A (Multiplier[6]), .B (p_0[6]), .CI (n_6));
FA_X1 i_6 (.CO (n_6), .S (p_1[5]), .A (Multiplier[5]), .B (p_0[5]), .CI (CLOCK_slo__sro_n1446));
INV_X1 slo__sro_c102 (.ZN (slo__sro_n163), .A (slo__n313));
FA_X1 i_4 (.CO (n_4), .S (p_1[3]), .A (Multiplier[3]), .B (p_0[3]), .CI (n_3));
FA_X1 i_3 (.CO (n_3), .S (p_1[2]), .A (Multiplier[2]), .B (p_0[2]), .CI (n_2));
FA_X1 i_2 (.CO (n_2), .S (p_1[1]), .A (Multiplier[1]), .B (p_0[1]), .CI (n_1));
HA_X1 i_1 (.CO (n_1), .S (p_1[0]), .A (Multiplier[0]), .B (p_0[0]));
XNOR2_X1 CLOCK_slo__sro_c975 (.ZN (CLOCK_slo__sro_n1249), .A (p_0[22]), .B (Multiplier[22]));
NOR2_X1 sgo__sro_c4 (.ZN (sgo__sro_n60), .A1 (n_33), .A2 (Multiplier[30]));
XNOR2_X1 CLOCK_slo__sro_c976 (.ZN (p_1[22]), .A (CLOCK_slo__sro_n1249), .B (n_22));
OR2_X1 sgo__sro_c6 (.ZN (sgo__sro_n58), .A1 (p_0[30]), .A2 (n_34));
OAI21_X2 sgo__sro_c7 (.ZN (sgo__sro_n57), .A (slo__mro_n810), .B1 (opt_ipo_n619), .B2 (sgo__sro_n58));
NAND2_X2 slo__sro_c30 (.ZN (slo__sro_n88), .A1 (p_0[29]), .A2 (Multiplier[29]));
NOR2_X4 slo__sro_c31 (.ZN (slo__sro_n87), .A1 (p_0[29]), .A2 (Multiplier[29]));
OAI21_X2 slo__sro_c32 (.ZN (slo__sro_n86), .A (slo__sro_n88), .B1 (slo__sro_n89), .B2 (slo__sro_n87));
XNOR2_X1 slo__sro_c33 (.ZN (slo__sro_n85), .A (p_0[29]), .B (Multiplier[29]));
XNOR2_X2 slo__sro_c34 (.ZN (p_1[29]), .A (slo__xsl_n846), .B (slo__sro_n85));
NAND2_X1 slo__sro_c51 (.ZN (slo__sro_n108), .A1 (p_0[4]), .A2 (Multiplier[4]));
NOR2_X2 slo__sro_c52 (.ZN (slo__sro_n107), .A1 (p_0[4]), .A2 (Multiplier[4]));
INV_X2 CLOCK_slo__sro_c1357 (.ZN (CLOCK_slo__sro_n1625), .A (slo__sro_n786));
XNOR2_X1 slo__sro_c54 (.ZN (slo__sro_n106), .A (p_0[4]), .B (Multiplier[4]));
XNOR2_X1 slo__sro_c55 (.ZN (p_1[4]), .A (slo__sro_n106), .B (n_4));
NAND2_X2 slo__sro_c103 (.ZN (slo__sro_n162), .A1 (slo__n353), .A2 (drc_ipoPP_0));
NOR2_X4 slo__sro_c104 (.ZN (slo__sro_n161), .A1 (slo__n353), .A2 (Multiplier[28]));
OAI21_X2 slo__sro_c105 (.ZN (slo__sro_n160), .A (slo__sro_n162), .B1 (slo__sro_n163), .B2 (slo__sro_n161));
XNOR2_X1 slo__sro_c106 (.ZN (slo__sro_n159), .A (p_0[28]), .B (Multiplier[28]));
XNOR2_X1 slo__sro_c107 (.ZN (p_1[28]), .A (n_28), .B (slo__sro_n159));
INV_X2 slo__sro_c77 (.ZN (slo__sro_n138), .A (n_14));
NAND2_X1 slo__sro_c78 (.ZN (slo__sro_n137), .A1 (p_0[14]), .A2 (Multiplier[14]));
NOR2_X1 slo__sro_c79 (.ZN (slo__sro_n136), .A1 (p_0[14]), .A2 (Multiplier[14]));
OAI21_X2 slo__sro_c80 (.ZN (slo__sro_n135), .A (slo__sro_n137), .B1 (slo__sro_n138), .B2 (slo__sro_n136));
XNOR2_X1 slo__sro_c81 (.ZN (slo__sro_n134), .A (p_0[14]), .B (Multiplier[14]));
XNOR2_X1 slo__sro_c82 (.ZN (p_1[14]), .A (slo__sro_n134), .B (n_14));
NOR2_X2 slo__sro_c122 (.ZN (slo__sro_n181), .A1 (p_0[27]), .A2 (Multiplier[27]));
OAI21_X1 slo__sro_c123 (.ZN (n_28), .A (slo__sro_n182), .B1 (slo__sro_n183), .B2 (slo__sro_n181));
XNOR2_X1 slo__sro_c124 (.ZN (slo__sro_n180), .A (p_0[27]), .B (Multiplier[27]));
XNOR2_X1 slo__sro_c125 (.ZN (p_1[27]), .A (slo__sro_n180), .B (n_27));
NAND2_X1 slo__sro_c144 (.ZN (slo__sro_n202), .A1 (p_0[19]), .A2 (Multiplier[19]));
NOR2_X1 slo__sro_c145 (.ZN (slo__sro_n201), .A1 (p_0[19]), .A2 (Multiplier[19]));
OAI21_X1 slo__sro_c146 (.ZN (slo__sro_n200), .A (slo__sro_n202), .B1 (slo__sro_n203), .B2 (slo__sro_n201));
XNOR2_X1 slo__sro_c147 (.ZN (slo__sro_n199), .A (p_0[19]), .B (Multiplier[19]));
XNOR2_X1 slo__sro_c148 (.ZN (p_1[19]), .A (slo__sro_n199), .B (n_19));
NAND2_X1 slo__sro_c161 (.ZN (slo__sro_n221), .A1 (p_0[18]), .A2 (Multiplier[18]));
NOR2_X1 slo__sro_c162 (.ZN (slo__sro_n220), .A1 (p_0[18]), .A2 (Multiplier[18]));
OAI21_X1 slo__sro_c163 (.ZN (n_19), .A (slo__sro_n221), .B1 (slo__sro_n222), .B2 (slo__sro_n220));
XNOR2_X1 slo__sro_c164 (.ZN (slo__sro_n219), .A (p_0[18]), .B (Multiplier[18]));
XNOR2_X1 slo__sro_c165 (.ZN (p_1[18]), .A (slo__sro_n219), .B (n_18));
NAND2_X1 slo__sro_c175 (.ZN (slo__sro_n235), .A1 (p_0[24]), .A2 (Multiplier[24]));
NOR2_X1 slo__sro_c176 (.ZN (slo__sro_n234), .A1 (p_0[24]), .A2 (Multiplier[24]));
OAI21_X2 slo__sro_c177 (.ZN (slo__sro_n233), .A (slo__sro_n235), .B1 (slo__sro_n236), .B2 (slo__sro_n234));
XNOR2_X1 slo__sro_c178 (.ZN (slo__sro_n232), .A (p_0[24]), .B (Multiplier[24]));
XNOR2_X1 slo__sro_c179 (.ZN (p_1[24]), .A (slo__sro_n232), .B (n_24));
NAND2_X1 slo__sro_c623 (.ZN (slo__sro_n771), .A1 (p_0[12]), .A2 (Multiplier[12]));
INV_X1 slo__sro_c471 (.ZN (slo__sro_n595), .A (p_0[13]));
OAI21_X1 slo__c234 (.ZN (slo__n313), .A (slo__sro_n182), .B1 (slo__sro_n183), .B2 (slo__sro_n181));
BUF_X4 slo__c259 (.Z (slo__n353), .A (p_0[28]));
INV_X2 slo__sro_c334 (.ZN (slo__sro_n456), .A (n_23));
INV_X1 slo__sro_c247 (.ZN (slo__sro_n328), .A (Multiplier[31]));
XNOR2_X2 slo__sro_c248 (.ZN (p_1[31]), .A (sgo__sro_n57), .B (slo__sro_n328));
NAND2_X1 slo__sro_c335 (.ZN (slo__sro_n455), .A1 (p_0[23]), .A2 (Multiplier[23]));
NOR2_X1 slo__sro_c336 (.ZN (slo__sro_n454), .A1 (p_0[23]), .A2 (Multiplier[23]));
OAI21_X1 slo__sro_c337 (.ZN (n_24), .A (slo__sro_n455), .B1 (slo__sro_n456), .B2 (slo__sro_n454));
XNOR2_X1 slo__sro_c338 (.ZN (slo__sro_n453), .A (p_0[23]), .B (Multiplier[23]));
XNOR2_X1 slo__sro_c339 (.ZN (p_1[23]), .A (slo__sro_n453), .B (CLOCK_slo__xsl_n1571));
INV_X1 slo__sro_c470 (.ZN (slo__sro_n596), .A (Multiplier[13]));
NAND2_X1 slo__sro_c472 (.ZN (slo__sro_n594), .A1 (p_0[13]), .A2 (Multiplier[13]));
NAND2_X1 slo__sro_c473 (.ZN (slo__sro_n593), .A1 (slo__sro_n595), .A2 (slo__sro_n596));
NAND2_X2 slo__sro_c474 (.ZN (slo__sro_n592), .A1 (slo__sro_n769), .A2 (slo__sro_n593));
NAND2_X2 slo__sro_c475 (.ZN (n_14), .A1 (slo__sro_n592), .A2 (slo__sro_n594));
XNOR2_X1 slo__sro_c476 (.ZN (slo__sro_n591), .A (p_0[13]), .B (Multiplier[13]));
XNOR2_X1 slo__sro_c477 (.ZN (p_1[13]), .A (slo__sro_n769), .B (slo__sro_n591));
OAI21_X2 slo__sro_c625 (.ZN (slo__sro_n769), .A (slo__sro_n771), .B1 (slo__sro_n772), .B2 (slo__sro_n770));
INV_X2 opt_ipo_c498 (.ZN (opt_ipo_n619), .A (slo__sro_n86));
NAND2_X1 slo__sro_c600 (.ZN (slo__sro_n736), .A1 (p_0[17]), .A2 (Multiplier[17]));
NOR2_X2 slo__sro_c601 (.ZN (slo__sro_n735), .A1 (p_0[17]), .A2 (Multiplier[17]));
OAI21_X2 slo__sro_c602 (.ZN (n_18), .A (slo__sro_n736), .B1 (slo__sro_n737), .B2 (slo__sro_n735));
XNOR2_X1 slo__sro_c603 (.ZN (slo__sro_n734), .A (p_0[17]), .B (Multiplier[17]));
XNOR2_X1 slo__sro_c604 (.ZN (p_1[17]), .A (n_17), .B (slo__sro_n734));
XNOR2_X1 slo__sro_c626 (.ZN (slo__sro_n768), .A (p_0[12]), .B (Multiplier[12]));
XNOR2_X1 slo__sro_c627 (.ZN (p_1[12]), .A (CLOCK_slo__xsl_n1478), .B (slo__sro_n768));
NAND2_X1 slo__sro_c637 (.ZN (slo__sro_n788), .A1 (p_0[25]), .A2 (Multiplier[25]));
NOR2_X2 slo__sro_c638 (.ZN (slo__sro_n787), .A1 (p_0[25]), .A2 (Multiplier[25]));
OAI21_X2 slo__sro_c639 (.ZN (slo__sro_n786), .A (slo__sro_n788), .B1 (slo__sro_n789), .B2 (slo__sro_n787));
XNOR2_X1 slo__sro_c640 (.ZN (slo__sro_n785), .A (p_0[25]), .B (Multiplier[25]));
XNOR2_X1 slo__sro_c641 (.ZN (p_1[25]), .A (slo__sro_n785), .B (slo__sro_n233));
OAI21_X2 CLOCK_slo__sro_c974 (.ZN (n_23), .A (CLOCK_slo__sro_n1251), .B1 (CLOCK_slo__sro_n1252), .B2 (CLOCK_slo__sro_n1250));
INV_X1 slo__xsl_c685 (.ZN (slo__xsl_n847), .A (slo__sro_n160));
OAI211_X1 slo__mro_c659 (.ZN (slo__mro_n810), .A (sgo__sro_n60), .B (slo__sro_n88)
    , .C1 (slo__sro_n89), .C2 (slo__sro_n87));
INV_X1 CLOCK_slo__sro_c971 (.ZN (CLOCK_slo__sro_n1252), .A (n_22));
NAND2_X1 CLOCK_slo__sro_c972 (.ZN (CLOCK_slo__sro_n1251), .A1 (p_0[22]), .A2 (Multiplier[22]));
NOR2_X1 CLOCK_slo__sro_c973 (.ZN (CLOCK_slo__sro_n1250), .A1 (p_0[22]), .A2 (Multiplier[22]));
NAND2_X1 CLOCK_slo__sro_c1048 (.ZN (CLOCK_slo__sro_n1317), .A1 (p_0[11]), .A2 (Multiplier[11]));
NOR2_X1 CLOCK_slo__sro_c1049 (.ZN (CLOCK_slo__sro_n1316), .A1 (p_0[11]), .A2 (Multiplier[11]));
OAI21_X2 CLOCK_slo__sro_c1050 (.ZN (n_12), .A (CLOCK_slo__sro_n1317), .B1 (CLOCK_slo__sro_n1318), .B2 (CLOCK_slo__sro_n1316));
XNOR2_X1 CLOCK_slo__sro_c1051 (.ZN (CLOCK_slo__sro_n1315), .A (p_0[11]), .B (Multiplier[11]));
XNOR2_X1 CLOCK_slo__sro_c1052 (.ZN (p_1[11]), .A (n_11), .B (CLOCK_slo__sro_n1315));
NAND2_X1 CLOCK_slo__sro_c1158 (.ZN (CLOCK_slo__sro_n1416), .A1 (p_0[15]), .A2 (Multiplier[15]));
NOR2_X1 CLOCK_slo__sro_c1159 (.ZN (CLOCK_slo__sro_n1415), .A1 (p_0[15]), .A2 (Multiplier[15]));
OAI21_X2 CLOCK_slo__sro_c1160 (.ZN (n_16), .A (CLOCK_slo__sro_n1416), .B1 (CLOCK_slo__sro_n1417), .B2 (CLOCK_slo__sro_n1415));
XNOR2_X1 CLOCK_slo__sro_c1161 (.ZN (CLOCK_slo__sro_n1414), .A (p_0[15]), .B (Multiplier[15]));
XNOR2_X1 CLOCK_slo__sro_c1162 (.ZN (p_1[15]), .A (CLOCK_slo__sro_n1414), .B (slo__sro_n135));
INV_X1 CLOCK_slo__xsl_c1302 (.ZN (CLOCK_slo__xsl_n1572), .A (n_23));
INV_X1 CLOCK_slo__xsl_c1303 (.ZN (CLOCK_slo__xsl_n1571), .A (CLOCK_slo__xsl_n1572));
NAND2_X1 CLOCK_slo__sro_c1358 (.ZN (CLOCK_slo__sro_n1624), .A1 (p_0[26]), .A2 (Multiplier[26]));
NOR2_X2 CLOCK_slo__sro_c1359 (.ZN (CLOCK_slo__sro_n1623), .A1 (p_0[26]), .A2 (Multiplier[26]));
INV_X1 CLOCK_slo__xsl_c1221 (.ZN (CLOCK_slo__xsl_n1479), .A (n_12));
INV_X1 CLOCK_slo__xsl_c1222 (.ZN (CLOCK_slo__xsl_n1478), .A (CLOCK_slo__xsl_n1479));
OAI21_X4 CLOCK_slo__sro_c1360 (.ZN (n_27), .A (CLOCK_slo__sro_n1624), .B1 (CLOCK_slo__sro_n1625), .B2 (CLOCK_slo__sro_n1623));
XNOR2_X1 CLOCK_slo__sro_c1361 (.ZN (CLOCK_slo__sro_n1622), .A (p_0[26]), .B (Multiplier[26]));
XNOR2_X1 CLOCK_slo__sro_c1362 (.ZN (p_1[26]), .A (CLOCK_slo__sro_n1622), .B (slo__sro_n786));

endmodule //datapath__0_246

module datapath__0_242 (opt_ipoPP_1, opt_ipoPP_11, p_0, p_1, p_2);

output [31:0] p_2;
input [31:0] p_0;
input [31:0] p_1;
input opt_ipoPP_1;
input opt_ipoPP_11;
wire slo__n1273;
wire CLOCK_slo__mro_n2064;
wire n_1;
wire n_2;
wire n_3;
wire n_4;
wire n_5;
wire n_6;
wire n_7;
wire n_8;
wire n_9;
wire n_10;
wire n_11;
wire slo__sro_n351;
wire n_15;
wire n_16;
wire n_17;
wire n_18;
wire slo__sro_n346;
wire n_20;
wire n_21;
wire n_22;
wire n_23;
wire n_24;
wire n_26;
wire n_27;
wire n_28;
wire n_29;
wire n_32;
wire n_0;
wire n_34;
wire n_33;
wire slo__sro_n65;
wire slo__sro_n66;
wire slo__sro_n67;
wire slo__sro_n68;
wire slo__sro_n69;
wire slo__sro_n89;
wire slo__sro_n90;
wire slo__sro_n91;
wire slo__sro_n1022;
wire slo__sro_n114;
wire slo__sro_n115;
wire slo__sro_n116;
wire slo__sro_n117;
wire slo__sro_n196;
wire slo__sro_n197;
wire slo__sro_n198;
wire slo__sro_n199;
wire slo__sro_n200;
wire slo__sro_n331;
wire slo__sro_n332;
wire slo__sro_n333;
wire slo__sro_n334;
wire slo__sro_n335;
wire slo__sro_n347;
wire slo__sro_n348;
wire slo__sro_n349;
wire slo__sro_n350;
wire slo__sro_n284;
wire slo__sro_n285;
wire slo__sro_n286;
wire slo__sro_n287;
wire slo__sro_n288;
wire slo__sro_n352;
wire slo__sro_n784;
wire slo__sro_n372;
wire slo__sro_n373;
wire slo__sro_n374;
wire slo__sro_n375;
wire slo__sro_n462;
wire slo__sro_n463;
wire CLOCK_slo__sro_n1840;
wire slo__sro_n439;
wire slo__sro_n440;
wire slo__sro_n441;
wire slo__sro_n464;
wire slo__sro_n785;
wire slo__sro_n786;
wire slo__sro_n787;
wire slo__sro_n788;
wire slo__sro_n789;
wire slo__sro_n803;
wire slo__sro_n804;
wire slo__sro_n805;
wire slo__sro_n806;
wire slo__sro_n980;
wire slo__sro_n981;
wire slo__sro_n982;
wire slo__sro_n983;
wire slo__sro_n1023;
wire slo__sro_n1024;
wire slo__sro_n1025;
wire slo__sro_n1076;
wire slo__sro_n1077;
wire slo__sro_n1078;
wire slo__sro_n1079;
wire slo__sro_n1080;
wire slo__sro_n1115;
wire slo__sro_n1116;
wire slo__sro_n1117;
wire slo__sro_n1118;
wire slo__sro_n1514;
wire CLOCK_slo__sro_n1816;
wire CLOCK_slo__sro_n1817;
wire CLOCK_slo__sro_n1818;
wire CLOCK_slo__mro_n1827;
wire CLOCK_slo__sro_n1841;
wire CLOCK_slo__sro_n1842;
wire CLOCK_slo__sro_n1843;
wire CLOCK_slo__xsl_n1862;
wire CLOCK_slo__xsl_n1863;
wire CLOCK_slo__sro_n1874;
wire CLOCK_slo__sro_n1875;
wire CLOCK_slo__sro_n1876;
wire CLOCK_slo__sro_n1877;
wire CLOCK_slo__sro_n1891;
wire CLOCK_slo__sro_n1892;
wire CLOCK_slo__sro_n1893;
wire CLOCK_slo__sro_n1894;
wire CLOCK_slo__sro_n1895;
wire CLOCK_slo__sro_n1896;
wire CLOCK_slo__sro_n1924;
wire CLOCK_slo__sro_n1925;
wire CLOCK_slo__sro_n1926;
wire CLOCK_slo__sro_n1927;


INV_X1 i_36 (.ZN (n_34), .A (p_0[30]));
INV_X1 i_35 (.ZN (n_33), .A (p_1[30]));
INV_X1 i_34 (.ZN (n_32), .A (slo__sro_n66));
INV_X1 slo__sro_c652 (.ZN (slo__sro_n789), .A (p_0[9]));
OAI21_X2 CLOCK_slo__sro_c1410 (.ZN (n_27), .A (CLOCK_slo__sro_n1842), .B1 (CLOCK_slo__sro_n1841), .B2 (CLOCK_slo__sro_n1843));
OAI22_X1 i_31 (.ZN (n_0), .A1 (n_34), .A2 (p_1[30]), .B1 (p_0[30]), .B2 (n_33));
XNOR2_X1 i_0 (.ZN (p_2[30]), .A (n_32), .B (n_0));
INV_X2 slo__sro_c23 (.ZN (slo__sro_n91), .A (n_28));
NAND2_X1 slo__sro_c821 (.ZN (slo__sro_n1024), .A1 (p_1[27]), .A2 (p_0[27]));
INV_X1 slo__sro_c859 (.ZN (slo__sro_n1080), .A (n_24));
INV_X1 CLOCK_slo__xsl_c1432 (.ZN (CLOCK_slo__xsl_n1863), .A (n_11));
FA_X1 i_26 (.CO (n_26), .S (p_2[25]), .A (p_0[25]), .B (p_1[25]), .CI (slo__sro_n1077));
INV_X1 slo__sro_c892 (.ZN (slo__sro_n1118), .A (n_7));
INV_X1 CLOCK_slo__sro_c1458 (.ZN (CLOCK_slo__sro_n1896), .A (p_0[22]));
INV_X1 CLOCK_slo__sro_c1491 (.ZN (CLOCK_slo__sro_n1927), .A (n_3));
FA_X1 i_22 (.CO (n_22), .S (p_2[21]), .A (p_0[21]), .B (p_1[21]), .CI (n_21));
FA_X1 i_21 (.CO (n_21), .S (p_2[20]), .A (p_0[20]), .B (p_1[20]), .CI (n_20));
FA_X1 i_20 (.CO (n_20), .S (p_2[19]), .A (p_0[19]), .B (p_1[19]), .CI (slo__sro_n332));
INV_X1 slo__sro_c264 (.ZN (slo__sro_n352), .A (n_34));
NAND2_X1 slo__sro_c654 (.ZN (slo__sro_n787), .A1 (p_1[9]), .A2 (p_0[9]));
NOR2_X1 slo__sro_c822 (.ZN (slo__sro_n1023), .A1 (p_1[27]), .A2 (p_0[27]));
XNOR2_X2 CLOCK_slo__mro_c1397 (.ZN (CLOCK_slo__mro_n1827), .A (n_10), .B (p_0[10]));
FA_X1 i_15 (.CO (n_15), .S (p_2[14]), .A (p_0[14]), .B (p_1[14]), .CI (slo__sro_n285));
INV_X1 slo__sro_c653 (.ZN (slo__sro_n788), .A (p_1[9]));
NAND2_X1 slo__sro_c365 (.ZN (slo__sro_n464), .A1 (p_1[17]), .A2 (p_0[17]));
INV_X2 slo__sro_c250 (.ZN (slo__sro_n335), .A (n_18));
XNOR2_X1 slo__sro_c368 (.ZN (slo__sro_n462), .A (p_1[17]), .B (p_0[17]));
INV_X1 slo__sro_c670 (.ZN (slo__sro_n806), .A (n_8));
INV_X2 slo__sro_c780 (.ZN (slo__sro_n983), .A (n_16));
OAI21_X2 slo__c1007 (.ZN (slo__n1273), .A (slo__sro_n982), .B1 (slo__sro_n983), .B2 (slo__sro_n981));
INV_X1 slo__sro_c129 (.ZN (slo__sro_n200), .A (n_11));
FA_X1 i_6 (.CO (n_6), .S (p_2[5]), .A (p_0[5]), .B (p_1[5]), .CI (n_5));
FA_X1 i_5 (.CO (n_5), .S (p_2[4]), .A (p_0[4]), .B (p_1[4]), .CI (n_4));
XNOR2_X1 CLOCK_slo__mro_c1593 (.ZN (CLOCK_slo__mro_n2064), .A (p_1[28]), .B (p_0[28]));
FA_X1 i_3 (.CO (n_3), .S (p_2[2]), .A (p_0[2]), .B (p_1[2]), .CI (n_2));
FA_X1 i_2 (.CO (n_2), .S (p_2[1]), .A (p_0[1]), .B (p_1[1]), .CI (n_1));
HA_X1 i_1 (.CO (n_1), .S (p_2[0]), .A (p_0[0]), .B (p_1[0]));
INV_X2 slo__sro_c3 (.ZN (slo__sro_n69), .A (n_29));
NAND2_X1 slo__sro_c4 (.ZN (slo__sro_n68), .A1 (p_1[29]), .A2 (p_0[29]));
NOR2_X1 slo__sro_c5 (.ZN (slo__sro_n67), .A1 (p_1[29]), .A2 (p_0[29]));
OAI21_X2 slo__sro_c6 (.ZN (slo__sro_n66), .A (slo__sro_n68), .B1 (slo__sro_n69), .B2 (slo__sro_n67));
XNOR2_X2 slo__sro_c7 (.ZN (slo__sro_n65), .A (p_1[29]), .B (p_0[29]));
XNOR2_X1 slo__sro_c8 (.ZN (p_2[29]), .A (n_29), .B (slo__sro_n65));
NAND2_X1 slo__sro_c24 (.ZN (slo__sro_n90), .A1 (p_1[28]), .A2 (p_0[28]));
NOR2_X1 slo__sro_c25 (.ZN (slo__sro_n89), .A1 (p_1[28]), .A2 (p_0[28]));
OAI21_X2 slo__sro_c26 (.ZN (n_29), .A (slo__sro_n90), .B1 (slo__sro_n89), .B2 (slo__sro_n91));
XNOR2_X1 slo__sro_c28 (.ZN (p_2[28]), .A (CLOCK_slo__mro_n2064), .B (n_28));
INV_X2 slo__sro_c820 (.ZN (slo__sro_n1025), .A (n_27));
INV_X1 slo__sro_c50 (.ZN (slo__sro_n117), .A (n_6));
NAND2_X1 slo__sro_c51 (.ZN (slo__sro_n116), .A1 (p_1[6]), .A2 (p_0[6]));
NOR2_X1 slo__sro_c52 (.ZN (slo__sro_n115), .A1 (p_1[6]), .A2 (p_0[6]));
OAI21_X1 slo__sro_c53 (.ZN (n_7), .A (slo__sro_n116), .B1 (slo__sro_n117), .B2 (slo__sro_n115));
XNOR2_X1 slo__sro_c54 (.ZN (slo__sro_n114), .A (p_1[6]), .B (p_0[6]));
XNOR2_X1 slo__sro_c55 (.ZN (p_2[6]), .A (n_6), .B (slo__sro_n114));
NAND2_X1 slo__sro_c130 (.ZN (slo__sro_n199), .A1 (p_1[11]), .A2 (p_0[11]));
NOR2_X1 slo__sro_c131 (.ZN (slo__sro_n198), .A1 (p_1[11]), .A2 (p_0[11]));
OAI21_X2 slo__sro_c132 (.ZN (slo__sro_n197), .A (slo__sro_n199), .B1 (slo__sro_n200), .B2 (slo__sro_n198));
XNOR2_X1 slo__sro_c133 (.ZN (slo__sro_n196), .A (p_1[11]), .B (p_0[11]));
XNOR2_X2 slo__sro_c134 (.ZN (p_2[11]), .A (slo__sro_n196), .B (CLOCK_slo__xsl_n1862));
NAND2_X1 slo__sro_c251 (.ZN (slo__sro_n334), .A1 (p_1[18]), .A2 (p_0[18]));
NOR2_X2 slo__sro_c252 (.ZN (slo__sro_n333), .A1 (p_1[18]), .A2 (p_0[18]));
OAI21_X1 slo__sro_c253 (.ZN (slo__sro_n332), .A (slo__sro_n334), .B1 (slo__sro_n335), .B2 (slo__sro_n333));
XNOR2_X1 slo__sro_c254 (.ZN (slo__sro_n331), .A (p_1[18]), .B (p_0[18]));
XNOR2_X1 slo__sro_c255 (.ZN (p_2[18]), .A (slo__sro_n331), .B (n_18));
INV_X1 slo__sro_c265 (.ZN (slo__sro_n351), .A (p_1[30]));
INV_X1 slo__sro_c266 (.ZN (slo__sro_n350), .A (slo__sro_n66));
NOR2_X1 slo__sro_c267 (.ZN (slo__sro_n349), .A1 (n_33), .A2 (p_0[30]));
NAND2_X1 slo__sro_c268 (.ZN (slo__sro_n348), .A1 (slo__sro_n349), .A2 (slo__sro_n350));
NAND2_X1 slo__sro_c269 (.ZN (slo__sro_n347), .A1 (slo__sro_n351), .A2 (slo__sro_n352));
OAI21_X2 slo__sro_c270 (.ZN (slo__sro_n346), .A (slo__sro_n348), .B1 (n_32), .B2 (slo__sro_n347));
INV_X1 slo__sro_c210 (.ZN (slo__sro_n288), .A (slo__sro_n373));
NAND2_X1 slo__sro_c211 (.ZN (slo__sro_n287), .A1 (p_1[13]), .A2 (p_0[13]));
NOR2_X1 slo__sro_c212 (.ZN (slo__sro_n286), .A1 (p_1[13]), .A2 (p_0[13]));
OAI21_X2 slo__sro_c213 (.ZN (slo__sro_n285), .A (slo__sro_n287), .B1 (slo__sro_n288), .B2 (slo__sro_n286));
XNOR2_X1 slo__sro_c214 (.ZN (slo__sro_n284), .A (opt_ipoPP_1), .B (p_0[13]));
XNOR2_X1 slo__sro_c215 (.ZN (p_2[13]), .A (slo__sro_n284), .B (slo__sro_n373));
NAND2_X1 slo__sro_c286 (.ZN (slo__sro_n375), .A1 (p_1[12]), .A2 (p_0[12]));
OAI21_X4 slo__sro_c287 (.ZN (slo__sro_n374), .A (slo__sro_n197), .B1 (p_1[12]), .B2 (p_0[12]));
NAND2_X4 slo__sro_c288 (.ZN (slo__sro_n373), .A1 (slo__sro_n374), .A2 (slo__sro_n375));
XNOR2_X1 slo__sro_c289 (.ZN (slo__sro_n372), .A (p_1[12]), .B (p_0[12]));
XNOR2_X1 slo__sro_c290 (.ZN (p_2[12]), .A (slo__sro_n372), .B (slo__sro_n197));
OAI21_X2 slo__sro_c366 (.ZN (slo__sro_n463), .A (slo__n1273), .B1 (p_1[17]), .B2 (p_0[17]));
NAND2_X2 slo__sro_c367 (.ZN (n_18), .A1 (slo__sro_n463), .A2 (slo__sro_n464));
INV_X1 slo__sro_c342 (.ZN (slo__sro_n441), .A (n_10));
NAND2_X1 slo__sro_c343 (.ZN (slo__sro_n440), .A1 (p_1[10]), .A2 (p_0[10]));
NOR2_X1 slo__sro_c344 (.ZN (slo__sro_n439), .A1 (p_1[10]), .A2 (p_0[10]));
OAI21_X1 slo__sro_c345 (.ZN (n_11), .A (slo__sro_n440), .B1 (slo__sro_n439), .B2 (slo__sro_n441));
INV_X1 CLOCK_slo__sro_c1407 (.ZN (CLOCK_slo__sro_n1843), .A (n_26));
NAND2_X1 CLOCK_slo__sro_c1408 (.ZN (CLOCK_slo__sro_n1842), .A1 (p_0[26]), .A2 (p_1[26]));
XNOR2_X1 slo__sro_c369 (.ZN (p_2[17]), .A (slo__sro_n462), .B (n_17));
NAND2_X1 slo__sro_c655 (.ZN (slo__sro_n786), .A1 (slo__sro_n788), .A2 (slo__sro_n789));
NAND2_X1 slo__sro_c656 (.ZN (slo__sro_n785), .A1 (n_9), .A2 (slo__sro_n786));
NAND2_X2 slo__sro_c657 (.ZN (n_10), .A1 (slo__sro_n785), .A2 (slo__sro_n787));
XNOR2_X1 slo__sro_c658 (.ZN (slo__sro_n784), .A (p_1[9]), .B (p_0[9]));
XNOR2_X1 slo__sro_c659 (.ZN (p_2[9]), .A (n_9), .B (slo__sro_n784));
NAND2_X1 slo__sro_c671 (.ZN (slo__sro_n805), .A1 (p_1[8]), .A2 (p_0[8]));
NOR2_X1 slo__sro_c672 (.ZN (slo__sro_n804), .A1 (p_1[8]), .A2 (p_0[8]));
OAI21_X1 slo__sro_c673 (.ZN (n_9), .A (slo__sro_n805), .B1 (slo__sro_n806), .B2 (slo__sro_n804));
XNOR2_X1 slo__sro_c674 (.ZN (slo__sro_n803), .A (p_1[8]), .B (p_0[8]));
XNOR2_X1 slo__sro_c675 (.ZN (p_2[8]), .A (slo__sro_n803), .B (n_8));
NAND2_X1 slo__sro_c781 (.ZN (slo__sro_n982), .A1 (p_1[16]), .A2 (p_0[16]));
NOR2_X2 slo__sro_c782 (.ZN (slo__sro_n981), .A1 (p_1[16]), .A2 (p_0[16]));
OAI21_X1 slo__sro_c783 (.ZN (n_17), .A (slo__sro_n982), .B1 (slo__sro_n983), .B2 (slo__sro_n981));
XNOR2_X1 slo__sro_c784 (.ZN (slo__sro_n980), .A (p_1[16]), .B (p_0[16]));
XNOR2_X1 slo__sro_c785 (.ZN (p_2[16]), .A (slo__sro_n980), .B (n_16));
OAI21_X4 slo__sro_c823 (.ZN (n_28), .A (slo__sro_n1024), .B1 (slo__sro_n1025), .B2 (slo__sro_n1023));
XNOR2_X1 slo__sro_c824 (.ZN (slo__sro_n1022), .A (p_1[27]), .B (p_0[27]));
XNOR2_X1 slo__sro_c825 (.ZN (p_2[27]), .A (slo__sro_n1022), .B (n_27));
NAND2_X1 slo__sro_c860 (.ZN (slo__sro_n1079), .A1 (p_0[24]), .A2 (p_1[24]));
NOR2_X1 slo__sro_c861 (.ZN (slo__sro_n1078), .A1 (p_1[24]), .A2 (p_0[24]));
OAI21_X1 slo__sro_c862 (.ZN (slo__sro_n1077), .A (slo__sro_n1079), .B1 (slo__sro_n1080), .B2 (slo__sro_n1078));
XNOR2_X1 slo__sro_c863 (.ZN (slo__sro_n1076), .A (p_1[24]), .B (p_0[24]));
XNOR2_X1 slo__sro_c864 (.ZN (p_2[24]), .A (n_24), .B (slo__sro_n1076));
NAND2_X1 slo__sro_c893 (.ZN (slo__sro_n1117), .A1 (opt_ipoPP_11), .A2 (p_0[7]));
NOR2_X1 slo__sro_c894 (.ZN (slo__sro_n1116), .A1 (opt_ipoPP_11), .A2 (p_0[7]));
OAI21_X2 slo__sro_c895 (.ZN (n_8), .A (slo__sro_n1117), .B1 (slo__sro_n1118), .B2 (slo__sro_n1116));
XNOR2_X1 slo__sro_c896 (.ZN (slo__sro_n1115), .A (p_1[7]), .B (p_0[7]));
XNOR2_X1 slo__sro_c897 (.ZN (p_2[7]), .A (slo__sro_n1115), .B (n_7));
INV_X1 slo__sro_c1188 (.ZN (slo__sro_n1514), .A (p_0[31]));
XNOR2_X2 slo__sro_c1189 (.ZN (p_2[31]), .A (slo__sro_n346), .B (slo__sro_n1514));
NAND2_X1 CLOCK_slo__sro_c1385 (.ZN (CLOCK_slo__sro_n1818), .A1 (n_15), .A2 (p_0[15]));
AOI22_X2 CLOCK_slo__sro_c1386 (.ZN (CLOCK_slo__sro_n1817), .A1 (n_15), .A2 (p_1[15])
    , .B1 (p_1[15]), .B2 (p_0[15]));
NAND2_X2 CLOCK_slo__sro_c1387 (.ZN (n_16), .A1 (CLOCK_slo__sro_n1817), .A2 (CLOCK_slo__sro_n1818));
XNOR2_X1 CLOCK_slo__sro_c1388 (.ZN (CLOCK_slo__sro_n1816), .A (p_1[15]), .B (p_0[15]));
XNOR2_X1 CLOCK_slo__sro_c1389 (.ZN (p_2[15]), .A (CLOCK_slo__sro_n1816), .B (n_15));
XNOR2_X2 CLOCK_slo__mro_c1398 (.ZN (p_2[10]), .A (CLOCK_slo__mro_n1827), .B (p_1[10]));
NOR2_X1 CLOCK_slo__sro_c1409 (.ZN (CLOCK_slo__sro_n1841), .A1 (p_1[26]), .A2 (p_0[26]));
XNOR2_X1 CLOCK_slo__sro_c1411 (.ZN (CLOCK_slo__sro_n1840), .A (p_1[26]), .B (p_0[26]));
XNOR2_X1 CLOCK_slo__sro_c1412 (.ZN (p_2[26]), .A (CLOCK_slo__sro_n1840), .B (n_26));
INV_X1 CLOCK_slo__xsl_c1433 (.ZN (CLOCK_slo__xsl_n1862), .A (CLOCK_slo__xsl_n1863));
INV_X1 CLOCK_slo__sro_c1442 (.ZN (CLOCK_slo__sro_n1877), .A (n_23));
NAND2_X1 CLOCK_slo__sro_c1443 (.ZN (CLOCK_slo__sro_n1876), .A1 (p_1[23]), .A2 (p_0[23]));
NOR2_X1 CLOCK_slo__sro_c1444 (.ZN (CLOCK_slo__sro_n1875), .A1 (p_1[23]), .A2 (p_0[23]));
OAI21_X1 CLOCK_slo__sro_c1445 (.ZN (n_24), .A (CLOCK_slo__sro_n1876), .B1 (CLOCK_slo__sro_n1877), .B2 (CLOCK_slo__sro_n1875));
XNOR2_X2 CLOCK_slo__sro_c1446 (.ZN (CLOCK_slo__sro_n1874), .A (p_1[23]), .B (p_0[23]));
XNOR2_X2 CLOCK_slo__sro_c1447 (.ZN (p_2[23]), .A (n_23), .B (CLOCK_slo__sro_n1874));
INV_X1 CLOCK_slo__sro_c1459 (.ZN (CLOCK_slo__sro_n1895), .A (p_1[22]));
NAND2_X1 CLOCK_slo__sro_c1460 (.ZN (CLOCK_slo__sro_n1894), .A1 (p_1[22]), .A2 (p_0[22]));
NAND2_X1 CLOCK_slo__sro_c1461 (.ZN (CLOCK_slo__sro_n1893), .A1 (CLOCK_slo__sro_n1895), .A2 (CLOCK_slo__sro_n1896));
NAND2_X2 CLOCK_slo__sro_c1462 (.ZN (CLOCK_slo__sro_n1892), .A1 (n_22), .A2 (CLOCK_slo__sro_n1893));
NAND2_X1 CLOCK_slo__sro_c1463 (.ZN (n_23), .A1 (CLOCK_slo__sro_n1892), .A2 (CLOCK_slo__sro_n1894));
XNOR2_X1 CLOCK_slo__sro_c1464 (.ZN (CLOCK_slo__sro_n1891), .A (p_1[22]), .B (p_0[22]));
XNOR2_X1 CLOCK_slo__sro_c1465 (.ZN (p_2[22]), .A (n_22), .B (CLOCK_slo__sro_n1891));
NAND2_X1 CLOCK_slo__sro_c1492 (.ZN (CLOCK_slo__sro_n1926), .A1 (p_1[3]), .A2 (p_0[3]));
NOR2_X1 CLOCK_slo__sro_c1493 (.ZN (CLOCK_slo__sro_n1925), .A1 (p_1[3]), .A2 (p_0[3]));
OAI21_X1 CLOCK_slo__sro_c1494 (.ZN (n_4), .A (CLOCK_slo__sro_n1926), .B1 (CLOCK_slo__sro_n1927), .B2 (CLOCK_slo__sro_n1925));
XNOR2_X2 CLOCK_slo__sro_c1495 (.ZN (CLOCK_slo__sro_n1924), .A (p_1[3]), .B (p_0[3]));
XNOR2_X1 CLOCK_slo__sro_c1496 (.ZN (p_2[3]), .A (CLOCK_slo__sro_n1924), .B (n_3));

endmodule //datapath__0_242

module datapath__0_241 (p_0_16_PP_0, p_0_16_PP_1, p_0_15_PP_0, Multiplier, p_0, p_1);

output [31:0] p_1;
input [31:0] Multiplier;
input [31:0] p_0;
input p_0_16_PP_0;
input p_0_16_PP_1;
input p_0_15_PP_0;
wire slo__n512;
wire slo_n532;
wire CLOCK_slo__sro_n1150;
wire n_1;
wire n_2;
wire n_3;
wire n_4;
wire n_5;
wire slo__sro_n477;
wire n_7;
wire n_8;
wire n_9;
wire n_10;
wire n_11;
wire n_13;
wire slo__sro_n257;
wire n_15;
wire n_16;
wire CLOCK_slo__sro_n1214;
wire n_19;
wire n_20;
wire n_23;
wire n_24;
wire n_25;
wire n_28;
wire n_30;
wire n_32;
wire n_0;
wire n_34;
wire n_33;
wire slo__sro_n63;
wire slo__sro_n64;
wire slo__sro_n65;
wire slo__sro_n66;
wire slo__sro_n100;
wire slo__sro_n101;
wire slo__sro_n102;
wire slo__sro_n103;
wire slo__sro_n128;
wire slo__sro_n129;
wire slo__sro_n130;
wire slo__sro_n131;
wire slo__sro_n132;
wire slo__sro_n148;
wire slo__sro_n149;
wire slo__sro_n150;
wire slo__sro_n151;
wire slo__sro_n191;
wire slo__sro_n192;
wire slo__sro_n193;
wire slo__sro_n194;
wire slo__sro_n195;
wire slo__sro_n208;
wire slo__sro_n209;
wire slo__sro_n210;
wire slo__sro_n211;
wire slo__sro_n212;
wire slo__sro_n225;
wire slo__sro_n226;
wire slo__sro_n227;
wire slo__sro_n228;
wire slo__sro_n229;
wire slo__sro_n242;
wire slo__sro_n243;
wire slo__sro_n244;
wire slo__sro_n245;
wire slo__sro_n246;
wire slo__sro_n258;
wire slo__sro_n259;
wire slo__sro_n476;
wire CLOCK_slo__sro_n1419;
wire slo__sro_n596;
wire slo__sro_n597;
wire CLOCK_slo__sro_n1418;
wire slo__sro_n378;
wire slo__sro_n379;
wire slo__sro_n380;
wire slo__sro_n381;
wire slo__sro_n478;
wire slo__sro_n479;
wire slo__sro_n481;
wire slo__sro_n598;
wire slo__sro_n599;
wire slo__sro_n647;
wire slo__sro_n648;
wire slo__sro_n649;
wire slo__sro_n650;
wire slo__sro_n651;
wire slo__mro_n677;
wire slo__sro_n751;
wire slo__sro_n752;
wire slo__sro_n753;
wire slo__sro_n754;
wire slo__sro_n755;
wire CLOCK_slo__sro_n1149;
wire slo__sro_n827;
wire slo__sro_n828;
wire slo__sro_n829;
wire CLOCK_slo__sro_n1080;
wire CLOCK_slo__sro_n1081;
wire CLOCK_slo__sro_n1082;
wire CLOCK_slo__sro_n1083;
wire CLOCK_slo__sro_n1110;
wire CLOCK_slo__n1446;
wire CLOCK_slo__sro_n1112;
wire CLOCK_slo__mro_n1125;
wire CLOCK_slo__sro_n1151;
wire CLOCK_slo__sro_n1152;
wire CLOCK_slo__sro_n1153;
wire CLOCK_slo__sro_n1154;
wire CLOCK_slo__mro_n1168;
wire CLOCK_slo__sro_n1215;
wire CLOCK_slo__sro_n1216;
wire CLOCK_slo__sro_n1217;
wire CLOCK_slo__mro_n1263;
wire CLOCK_slo__sro_n1420;
wire CLOCK_slo__sro_n1421;
wire CLOCK_slo__sro_n1451;
wire CLOCK_slo__sro_n1452;
wire CLOCK_slo__sro_n1453;
wire CLOCK_slo__sro_n1454;


INV_X1 i_36 (.ZN (n_34), .A (Multiplier[30]));
INV_X2 i_35 (.ZN (n_33), .A (p_0[30]));
INV_X4 i_34 (.ZN (n_32), .A (n_30));
INV_X1 slo__L4_c4_c380 (.ZN (slo_n532), .A (slo__n512));
NAND2_X1 slo__sro_c535 (.ZN (slo__sro_n754), .A1 (p_0[11]), .A2 (Multiplier[11]));
OAI22_X1 i_31 (.ZN (n_0), .A1 (n_34), .A2 (p_0[30]), .B1 (n_33), .B2 (Multiplier[30]));
XNOR2_X2 i_0 (.ZN (p_1[30]), .A (n_0), .B (n_32));
INV_X1 slo__sro_c47 (.ZN (slo__sro_n103), .A (slo__sro_n378));
INV_X2 slo__sro_c132 (.ZN (slo__sro_n195), .A (slo__sro_n129));
INV_X1 CLOCK_slo__sro_c817 (.ZN (CLOCK_slo__sro_n1154), .A (Multiplier[19]));
XNOR2_X1 slo__sro_c643 (.ZN (p_1[11]), .A (n_11), .B (slo__sro_n751));
INV_X1 slo__sro_c174 (.ZN (slo__sro_n246), .A (n_13));
FA_X1 i_25 (.CO (n_25), .S (p_1[24]), .A (Multiplier[24]), .B (p_0[24]), .CI (n_24));
FA_X1 i_24 (.CO (n_24), .S (p_1[23]), .A (Multiplier[23]), .B (p_0[23]), .CI (n_23));
FA_X1 i_23 (.CO (n_23), .S (p_1[22]), .A (Multiplier[22]), .B (p_0[22]), .CI (slo__sro_n209));
INV_X1 slo__sro_c160 (.ZN (slo__sro_n229), .A (n_25));
INV_X1 slo__mro_c477 (.ZN (slo__mro_n677), .A (Multiplier[31]));
XNOR2_X2 CLOCK_slo__mro_c837 (.ZN (CLOCK_slo__mro_n1168), .A (p_0[28]), .B (Multiplier[28]));
FA_X1 i_19 (.CO (n_19), .S (p_1[18]), .A (Multiplier[18]), .B (p_0[18]), .CI (slo__sro_n192));
INV_X1 slo__sro_c146 (.ZN (slo__sro_n212), .A (slo__sro_n648));
INV_X2 slo__sro_c90 (.ZN (slo__sro_n151), .A (n_28));
XNOR2_X2 slo__sro_c430 (.ZN (slo__sro_n596), .A (p_0[12]), .B (Multiplier[12]));
FA_X1 i_15 (.CO (n_15), .S (p_1[14]), .A (Multiplier[14]), .B (p_0[14]), .CI (slo__sro_n243));
OR2_X2 slo__sro_c188 (.ZN (slo__sro_n259), .A1 (n_33), .A2 (Multiplier[30]));
INV_X2 slo__sro_c452 (.ZN (slo__sro_n651), .A (n_20));
NAND2_X1 slo__sro_c596 (.ZN (slo__sro_n829), .A1 (p_0[26]), .A2 (Multiplier[26]));
OAI22_X2 CLOCK_slo__mro_c912 (.ZN (slo__sro_n257), .A1 (n_32), .A2 (slo__sro_n258)
    , .B1 (slo__sro_n259), .B2 (n_30));
FA_X1 i_10 (.CO (n_10), .S (p_1[9]), .A (Multiplier[9]), .B (p_0[9]), .CI (n_9));
FA_X1 i_9 (.CO (n_9), .S (p_1[8]), .A (Multiplier[8]), .B (p_0[8]), .CI (n_8));
FA_X1 i_8 (.CO (n_8), .S (p_1[7]), .A (Multiplier[7]), .B (p_0[7]), .CI (n_7));
INV_X2 slo__sro_c74 (.ZN (slo__sro_n132), .A (n_16));
NAND2_X1 slo__sro_c351 (.ZN (slo__sro_n479), .A1 (slo_n532), .A2 (Multiplier[15]));
FA_X1 i_4 (.CO (n_4), .S (p_1[3]), .A (Multiplier[3]), .B (p_0[3]), .CI (n_3));
FA_X1 i_2 (.CO (n_2), .S (p_1[1]), .A (Multiplier[1]), .B (p_0[1]), .CI (n_1));
HA_X1 i_1 (.CO (n_1), .S (p_1[0]), .A (Multiplier[0]), .B (p_0[0]));
INV_X2 slo__sro_c7 (.ZN (slo__sro_n66), .A (slo__sro_n148));
NAND2_X1 slo__sro_c8 (.ZN (slo__sro_n65), .A1 (p_0[29]), .A2 (Multiplier[29]));
NOR2_X2 slo__sro_c9 (.ZN (slo__sro_n64), .A1 (p_0[29]), .A2 (Multiplier[29]));
OAI21_X4 slo__sro_c10 (.ZN (n_30), .A (slo__sro_n65), .B1 (slo__sro_n66), .B2 (slo__sro_n64));
XNOR2_X2 slo__sro_c11 (.ZN (slo__sro_n63), .A (p_0[29]), .B (Multiplier[29]));
XNOR2_X2 slo__sro_c12 (.ZN (p_1[29]), .A (slo__sro_n63), .B (slo__sro_n148));
NAND2_X1 slo__sro_c48 (.ZN (slo__sro_n102), .A1 (p_0[6]), .A2 (Multiplier[6]));
NOR2_X1 slo__sro_c49 (.ZN (slo__sro_n101), .A1 (p_0[6]), .A2 (Multiplier[6]));
OAI21_X1 slo__sro_c50 (.ZN (n_7), .A (slo__sro_n102), .B1 (slo__sro_n101), .B2 (slo__sro_n103));
XNOR2_X1 slo__sro_c51 (.ZN (slo__sro_n100), .A (p_0[6]), .B (Multiplier[6]));
XNOR2_X1 slo__sro_c52 (.ZN (p_1[6]), .A (slo__sro_n100), .B (slo__sro_n378));
NAND2_X1 slo__sro_c75 (.ZN (slo__sro_n131), .A1 (p_0[16]), .A2 (Multiplier[16]));
NOR2_X1 slo__sro_c76 (.ZN (slo__sro_n130), .A1 (p_0_16_PP_0), .A2 (Multiplier[16]));
OAI21_X2 slo__sro_c77 (.ZN (slo__sro_n129), .A (slo__sro_n131), .B1 (slo__sro_n132), .B2 (slo__sro_n130));
XNOR2_X1 slo__sro_c78 (.ZN (slo__sro_n128), .A (p_0_16_PP_1), .B (Multiplier[16]));
XNOR2_X1 slo__sro_c79 (.ZN (p_1[16]), .A (slo__sro_n128), .B (n_16));
NAND2_X1 slo__sro_c91 (.ZN (slo__sro_n150), .A1 (p_0[28]), .A2 (Multiplier[28]));
NOR2_X1 slo__sro_c92 (.ZN (slo__sro_n149), .A1 (p_0[28]), .A2 (Multiplier[28]));
OAI21_X2 slo__sro_c93 (.ZN (slo__sro_n148), .A (slo__sro_n150), .B1 (slo__sro_n149), .B2 (slo__sro_n151));
INV_X1 CLOCK_slo__sro_c878 (.ZN (CLOCK_slo__sro_n1217), .A (n_10));
NAND2_X1 CLOCK_slo__sro_c879 (.ZN (CLOCK_slo__sro_n1216), .A1 (p_0[10]), .A2 (Multiplier[10]));
NAND2_X1 slo__sro_c133 (.ZN (slo__sro_n194), .A1 (p_0[17]), .A2 (Multiplier[17]));
NOR2_X1 slo__sro_c134 (.ZN (slo__sro_n193), .A1 (p_0[17]), .A2 (Multiplier[17]));
OAI21_X2 slo__sro_c135 (.ZN (slo__sro_n192), .A (slo__sro_n194), .B1 (slo__sro_n195), .B2 (slo__sro_n193));
XNOR2_X1 slo__sro_c136 (.ZN (slo__sro_n191), .A (p_0[17]), .B (Multiplier[17]));
XNOR2_X1 slo__sro_c137 (.ZN (p_1[17]), .A (slo__sro_n191), .B (slo__sro_n129));
NAND2_X1 slo__sro_c147 (.ZN (slo__sro_n211), .A1 (p_0[21]), .A2 (Multiplier[21]));
NOR2_X2 slo__sro_c148 (.ZN (slo__sro_n210), .A1 (p_0[21]), .A2 (Multiplier[21]));
OAI21_X1 slo__sro_c149 (.ZN (slo__sro_n209), .A (slo__sro_n211), .B1 (slo__sro_n212), .B2 (slo__sro_n210));
XNOR2_X1 slo__sro_c150 (.ZN (slo__sro_n208), .A (p_0[21]), .B (Multiplier[21]));
XNOR2_X1 slo__sro_c151 (.ZN (p_1[21]), .A (slo__sro_n208), .B (slo__sro_n648));
NAND2_X1 slo__sro_c161 (.ZN (slo__sro_n228), .A1 (p_0[25]), .A2 (Multiplier[25]));
NOR2_X2 slo__sro_c162 (.ZN (slo__sro_n227), .A1 (p_0[25]), .A2 (Multiplier[25]));
OAI21_X2 slo__sro_c163 (.ZN (slo__sro_n226), .A (slo__sro_n228), .B1 (slo__sro_n229), .B2 (slo__sro_n227));
XNOR2_X2 slo__sro_c164 (.ZN (slo__sro_n225), .A (p_0[25]), .B (Multiplier[25]));
XNOR2_X1 slo__sro_c165 (.ZN (p_1[25]), .A (slo__sro_n225), .B (n_25));
NAND2_X1 slo__sro_c175 (.ZN (slo__sro_n245), .A1 (p_0[13]), .A2 (Multiplier[13]));
NOR2_X1 slo__sro_c176 (.ZN (slo__sro_n244), .A1 (p_0[13]), .A2 (Multiplier[13]));
OAI21_X1 slo__sro_c177 (.ZN (slo__sro_n243), .A (slo__sro_n245), .B1 (slo__sro_n246), .B2 (slo__sro_n244));
XNOR2_X1 slo__sro_c178 (.ZN (slo__sro_n242), .A (p_0[13]), .B (Multiplier[13]));
XNOR2_X1 slo__sro_c179 (.ZN (p_1[13]), .A (n_13), .B (slo__sro_n242));
INV_X1 CLOCK_slo__sro_c1110 (.ZN (CLOCK_slo__sro_n1454), .A (n_2));
INV_X1 slo__sro_c534 (.ZN (slo__sro_n755), .A (n_11));
INV_X1 slo__L3_c3_c381 (.ZN (slo__n512), .A (p_0_15_PP_0));
NAND2_X1 slo__sro_c427 (.ZN (slo__sro_n598), .A1 (Multiplier[12]), .A2 (p_0[12]));
INV_X1 slo__sro_c349 (.ZN (slo__sro_n481), .A (Multiplier[15]));
INV_X1 slo__sro_c426 (.ZN (slo__sro_n599), .A (slo__sro_n752));
INV_X1 slo__sro_c266 (.ZN (slo__sro_n381), .A (n_5));
OAI21_X2 slo__sro_c429 (.ZN (n_13), .A (slo__sro_n598), .B1 (slo__sro_n599), .B2 (slo__sro_n597));
NOR2_X1 slo__sro_c428 (.ZN (slo__sro_n597), .A1 (p_0[12]), .A2 (Multiplier[12]));
NAND2_X1 slo__sro_c267 (.ZN (slo__sro_n380), .A1 (p_0[5]), .A2 (Multiplier[5]));
NOR2_X1 slo__sro_c268 (.ZN (slo__sro_n379), .A1 (p_0[5]), .A2 (Multiplier[5]));
OAI21_X1 slo__sro_c269 (.ZN (slo__sro_n378), .A (slo__sro_n380), .B1 (slo__sro_n381), .B2 (slo__sro_n379));
NOR2_X1 CLOCK_slo__c1101 (.ZN (CLOCK_slo__n1446), .A1 (p_0[30]), .A2 (n_34));
INV_X1 CLOCK_slo__sro_c1066 (.ZN (CLOCK_slo__sro_n1421), .A (p_0[27]));
NAND2_X1 slo__sro_c352 (.ZN (slo__sro_n478), .A1 (slo__n512), .A2 (slo__sro_n481));
NAND2_X1 slo__sro_c353 (.ZN (slo__sro_n477), .A1 (n_15), .A2 (slo__sro_n478));
NAND2_X2 slo__sro_c354 (.ZN (n_16), .A1 (slo__sro_n477), .A2 (slo__sro_n479));
XNOR2_X1 slo__sro_c355 (.ZN (slo__sro_n476), .A (p_0[15]), .B (Multiplier[15]));
XNOR2_X1 slo__sro_c356 (.ZN (p_1[15]), .A (n_15), .B (slo__sro_n476));
XNOR2_X1 slo__sro_c431 (.ZN (p_1[12]), .A (slo__sro_n752), .B (slo__sro_n596));
NAND2_X1 slo__sro_c453 (.ZN (slo__sro_n650), .A1 (p_0[20]), .A2 (Multiplier[20]));
NOR2_X2 slo__sro_c454 (.ZN (slo__sro_n649), .A1 (p_0[20]), .A2 (Multiplier[20]));
OAI21_X2 slo__sro_c455 (.ZN (slo__sro_n648), .A (slo__sro_n650), .B1 (slo__sro_n651), .B2 (slo__sro_n649));
XNOR2_X1 slo__sro_c456 (.ZN (slo__sro_n647), .A (p_0[20]), .B (Multiplier[20]));
XNOR2_X1 slo__sro_c457 (.ZN (p_1[20]), .A (n_20), .B (slo__sro_n647));
XNOR2_X1 CLOCK_slo__mro_c933 (.ZN (CLOCK_slo__mro_n1263), .A (n_5), .B (Multiplier[5]));
XNOR2_X1 CLOCK_slo__mro_c934 (.ZN (p_1[5]), .A (CLOCK_slo__mro_n1263), .B (p_0[5]));
NOR2_X1 slo__sro_c536 (.ZN (slo__sro_n753), .A1 (p_0[11]), .A2 (Multiplier[11]));
OAI21_X1 slo__sro_c537 (.ZN (slo__sro_n752), .A (slo__sro_n754), .B1 (slo__sro_n755), .B2 (slo__sro_n753));
XNOR2_X1 slo__sro_c538 (.ZN (slo__sro_n751), .A (p_0[11]), .B (Multiplier[11]));
OAI21_X1 slo__sro_c597 (.ZN (slo__sro_n828), .A (slo__sro_n226), .B1 (p_0[26]), .B2 (Multiplier[26]));
NAND2_X2 slo__sro_c598 (.ZN (slo__sro_n827), .A1 (slo__sro_n828), .A2 (slo__sro_n829));
INV_X1 CLOCK_slo__sro_c818 (.ZN (CLOCK_slo__sro_n1153), .A (p_0[19]));
NAND2_X1 CLOCK_slo__sro_c819 (.ZN (CLOCK_slo__sro_n1152), .A1 (p_0[19]), .A2 (Multiplier[19]));
INV_X1 CLOCK_slo__sro_c745 (.ZN (CLOCK_slo__sro_n1083), .A (n_4));
NAND2_X1 CLOCK_slo__sro_c746 (.ZN (CLOCK_slo__sro_n1082), .A1 (p_0[4]), .A2 (Multiplier[4]));
NOR2_X1 CLOCK_slo__sro_c747 (.ZN (CLOCK_slo__sro_n1081), .A1 (p_0[4]), .A2 (Multiplier[4]));
OAI21_X1 CLOCK_slo__sro_c748 (.ZN (n_5), .A (CLOCK_slo__sro_n1082), .B1 (CLOCK_slo__sro_n1083), .B2 (CLOCK_slo__sro_n1081));
XNOR2_X1 CLOCK_slo__sro_c749 (.ZN (CLOCK_slo__sro_n1080), .A (p_0[4]), .B (Multiplier[4]));
XNOR2_X2 CLOCK_slo__sro_c750 (.ZN (p_1[4]), .A (CLOCK_slo__sro_n1080), .B (n_4));
NAND2_X1 CLOCK_slo__sro_c779 (.ZN (CLOCK_slo__sro_n1112), .A1 (p_0[27]), .A2 (Multiplier[27]));
INV_X1 CLOCK_slo__c1103 (.ZN (slo__sro_n258), .A (CLOCK_slo__n1446));
NAND2_X4 CLOCK_slo__sro_c781 (.ZN (n_28), .A1 (CLOCK_slo__sro_n1418), .A2 (CLOCK_slo__sro_n1112));
XNOR2_X1 CLOCK_slo__sro_c782 (.ZN (CLOCK_slo__sro_n1110), .A (p_0[27]), .B (Multiplier[27]));
XNOR2_X1 CLOCK_slo__sro_c783 (.ZN (p_1[27]), .A (CLOCK_slo__sro_n1110), .B (slo__sro_n827));
XNOR2_X2 CLOCK_slo__mro_c796 (.ZN (CLOCK_slo__mro_n1125), .A (p_0[26]), .B (Multiplier[26]));
XNOR2_X1 CLOCK_slo__mro_c797 (.ZN (p_1[26]), .A (CLOCK_slo__mro_n1125), .B (slo__sro_n226));
NAND2_X1 CLOCK_slo__sro_c820 (.ZN (CLOCK_slo__sro_n1151), .A1 (CLOCK_slo__sro_n1153), .A2 (CLOCK_slo__sro_n1154));
NAND2_X2 CLOCK_slo__sro_c821 (.ZN (CLOCK_slo__sro_n1150), .A1 (n_19), .A2 (CLOCK_slo__sro_n1151));
NAND2_X2 CLOCK_slo__sro_c822 (.ZN (n_20), .A1 (CLOCK_slo__sro_n1150), .A2 (CLOCK_slo__sro_n1152));
XNOR2_X1 CLOCK_slo__sro_c823 (.ZN (CLOCK_slo__sro_n1149), .A (p_0[19]), .B (Multiplier[19]));
XNOR2_X1 CLOCK_slo__sro_c824 (.ZN (p_1[19]), .A (CLOCK_slo__sro_n1149), .B (n_19));
XNOR2_X2 CLOCK_slo__mro_c838 (.ZN (p_1[28]), .A (CLOCK_slo__mro_n1168), .B (n_28));
NOR2_X1 CLOCK_slo__sro_c880 (.ZN (CLOCK_slo__sro_n1215), .A1 (p_0[10]), .A2 (Multiplier[10]));
OAI21_X1 CLOCK_slo__sro_c881 (.ZN (n_11), .A (CLOCK_slo__sro_n1216), .B1 (CLOCK_slo__sro_n1217), .B2 (CLOCK_slo__sro_n1215));
XNOR2_X1 CLOCK_slo__sro_c882 (.ZN (CLOCK_slo__sro_n1214), .A (p_0[10]), .B (Multiplier[10]));
XNOR2_X1 CLOCK_slo__sro_c883 (.ZN (p_1[10]), .A (n_10), .B (CLOCK_slo__sro_n1214));
XNOR2_X2 CLOCK_slo__mro_c913 (.ZN (p_1[31]), .A (slo__sro_n257), .B (slo__mro_n677));
INV_X1 CLOCK_slo__sro_c1067 (.ZN (CLOCK_slo__sro_n1420), .A (Multiplier[27]));
NAND2_X1 CLOCK_slo__sro_c1068 (.ZN (CLOCK_slo__sro_n1419), .A1 (CLOCK_slo__sro_n1421), .A2 (CLOCK_slo__sro_n1420));
NAND2_X2 CLOCK_slo__sro_c1069 (.ZN (CLOCK_slo__sro_n1418), .A1 (CLOCK_slo__sro_n1419), .A2 (slo__sro_n827));
NAND2_X1 CLOCK_slo__sro_c1111 (.ZN (CLOCK_slo__sro_n1453), .A1 (p_0[2]), .A2 (Multiplier[2]));
NOR2_X1 CLOCK_slo__sro_c1112 (.ZN (CLOCK_slo__sro_n1452), .A1 (p_0[2]), .A2 (Multiplier[2]));
OAI21_X1 CLOCK_slo__sro_c1113 (.ZN (n_3), .A (CLOCK_slo__sro_n1453), .B1 (CLOCK_slo__sro_n1454), .B2 (CLOCK_slo__sro_n1452));
XNOR2_X1 CLOCK_slo__sro_c1114 (.ZN (CLOCK_slo__sro_n1451), .A (p_0[2]), .B (Multiplier[2]));
XNOR2_X2 CLOCK_slo__sro_c1115 (.ZN (p_1[2]), .A (CLOCK_slo__sro_n1451), .B (n_2));

endmodule //datapath__0_241

module datapath__0_237 (p_0, p_1, p_2);

output [31:0] p_2;
input [31:0] p_0;
input [31:0] p_1;
wire slo__sro_n548;
wire slo__sro_n310;
wire slo__sro_n454;
wire CLOCK_slo__n1670;
wire n_1;
wire n_2;
wire n_3;
wire n_4;
wire n_5;
wire n_6;
wire n_7;
wire n_8;
wire n_9;
wire n_10;
wire n_12;
wire n_13;
wire n_14;
wire n_16;
wire n_17;
wire n_18;
wire n_19;
wire n_20;
wire n_22;
wire n_24;
wire n_25;
wire n_26;
wire n_27;
wire n_28;
wire n_29;
wire n_32;
wire n_0;
wire n_34;
wire n_33;
wire slo__sro_n67;
wire slo__sro_n68;
wire slo__sro_n69;
wire slo__sro_n70;
wire slo__sro_n71;
wire slo__sro_n108;
wire slo__sro_n109;
wire slo__sro_n110;
wire slo__sro_n111;
wire slo__sro_n121;
wire slo__sro_n122;
wire slo__sro_n123;
wire slo__sro_n124;
wire slo__sro_n149;
wire slo__sro_n150;
wire slo__sro_n151;
wire slo__sro_n152;
wire slo__sro_n177;
wire slo__sro_n178;
wire slo__sro_n179;
wire slo__sro_n180;
wire slo__sro_n194;
wire slo__sro_n195;
wire slo__sro_n196;
wire slo__sro_n197;
wire slo__sro_n198;
wire slo__sro_n266;
wire slo__sro_n267;
wire slo__sro_n268;
wire slo__sro_n269;
wire slo__sro_n270;
wire slo__sro_n283;
wire slo__sro_n284;
wire slo__sro_n285;
wire slo__sro_n286;
wire slo__sro_n287;
wire slo__sro_n311;
wire slo__sro_n312;
wire slo__sro_n313;
wire slo__sro_n314;
wire slo__sro_n315;
wire slo__sro_n453;
wire slo__sro_n432;
wire slo__sro_n433;
wire slo__sro_n434;
wire slo__sro_n435;
wire slo__sro_n436;
wire slo__sro_n455;
wire slo__sro_n456;
wire slo__sro_n549;
wire slo__sro_n550;
wire slo__sro_n551;
wire slo__sro_n751;
wire slo__sro_n752;
wire slo__sro_n753;
wire slo__sro_n754;
wire CLOCK_slo__sro_n1482;
wire CLOCK_slo__sro_n1454;
wire CLOCK_slo__sro_n1429;
wire CLOCK_slo__sro_n1430;
wire CLOCK_slo__sro_n1431;
wire CLOCK_slo__sro_n1432;
wire CLOCK_slo__sro_n1455;
wire CLOCK_slo__sro_n1456;
wire CLOCK_slo__sro_n1457;
wire CLOCK_slo__sro_n1483;
wire CLOCK_slo__sro_n1484;
wire CLOCK_slo__sro_n1485;
wire CLOCK_slo__sro_n1486;
wire CLOCK_slo__sro_n1487;
wire CLOCK_slo__sro_n1623;
wire CLOCK_slo__sro_n1624;
wire CLOCK_slo__sro_n1625;


INV_X1 i_36 (.ZN (n_34), .A (p_0[30]));
INV_X1 i_35 (.ZN (n_33), .A (p_1[30]));
INV_X1 i_34 (.ZN (n_32), .A (slo__sro_n68));
NAND2_X1 slo__sro_c334 (.ZN (slo__sro_n455), .A1 (p_1[28]), .A2 (p_0[28]));
XOR2_X2 i_32 (.Z (p_2[31]), .A (slo__sro_n310), .B (p_0[31]));
OAI22_X1 i_31 (.ZN (n_0), .A1 (n_34), .A2 (p_1[30]), .B1 (n_33), .B2 (p_0[30]));
XNOR2_X1 i_0 (.ZN (p_2[30]), .A (n_32), .B (n_0));
INV_X1 slo__sro_c45 (.ZN (slo__sro_n111), .A (CLOCK_slo__n1670));
NAND2_X1 slo__sro_c415 (.ZN (slo__sro_n550), .A1 (p_1[16]), .A2 (p_0[16]));
NAND2_X1 CLOCK_slo__sro_c985 (.ZN (CLOCK_slo__sro_n1485), .A1 (p_1[8]), .A2 (p_0[8]));
FA_X1 i_27 (.CO (n_27), .S (p_2[26]), .A (p_0[26]), .B (p_1[26]), .CI (n_26));
FA_X1 i_26 (.CO (n_26), .S (p_2[25]), .A (p_0[25]), .B (p_1[25]), .CI (n_25));
INV_X2 slo__sro_c131 (.ZN (slo__sro_n198), .A (n_14));
INV_X1 slo__sro_c243 (.ZN (slo__sro_n315), .A (slo__sro_n68));
FA_X1 i_22 (.CO (n_22), .S (p_2[21]), .A (p_0[21]), .B (p_1[21]), .CI (slo__sro_n433));
OAI21_X2 slo__sro_c336 (.ZN (n_29), .A (slo__sro_n455), .B1 (slo__sro_n456), .B2 (slo__sro_n454));
XNOR2_X1 CLOCK_slo__sro_c929 (.ZN (p_2[9]), .A (CLOCK_slo__sro_n1429), .B (n_9));
FA_X1 i_19 (.CO (n_19), .S (p_2[18]), .A (p_0[18]), .B (p_1[18]), .CI (n_18));
INV_X2 slo__sro_c59 (.ZN (slo__sro_n124), .A (slo__sro_n195));
INV_X1 slo__sro_c86 (.ZN (slo__sro_n152), .A (n_7));
INV_X1 slo__sro_c207 (.ZN (slo__sro_n270), .A (n_10));
FA_X1 i_14 (.CO (n_14), .S (p_2[13]), .A (p_0[13]), .B (p_1[13]), .CI (n_13));
FA_X1 i_13 (.CO (n_13), .S (p_2[12]), .A (p_0[12]), .B (p_1[12]), .CI (n_12));
FA_X1 i_12 (.CO (n_12), .S (p_2[11]), .A (p_0[11]), .B (p_1[11]), .CI (slo__sro_n267));
INV_X1 slo__sro_c221 (.ZN (slo__sro_n287), .A (n_22));
INV_X1 CLOCK_slo__sro_c983 (.ZN (CLOCK_slo__sro_n1487), .A (p_0[8]));
NAND2_X1 slo__sro_c113 (.ZN (slo__sro_n180), .A1 (p_1[24]), .A2 (p_0[24]));
FA_X1 i_7 (.CO (n_7), .S (p_2[6]), .A (p_0[6]), .B (p_1[6]), .CI (n_6));
FA_X1 i_6 (.CO (n_6), .S (p_2[5]), .A (p_0[5]), .B (p_1[5]), .CI (n_5));
FA_X1 i_5 (.CO (n_5), .S (p_2[4]), .A (p_0[4]), .B (p_1[4]), .CI (n_4));
FA_X1 i_4 (.CO (n_4), .S (p_2[3]), .A (p_0[3]), .B (p_1[3]), .CI (n_3));
FA_X1 i_3 (.CO (n_3), .S (p_2[2]), .A (p_0[2]), .B (p_1[2]), .CI (n_2));
FA_X1 i_2 (.CO (n_2), .S (p_2[1]), .A (p_0[1]), .B (p_1[1]), .CI (n_1));
HA_X1 i_1 (.CO (n_1), .S (p_2[0]), .A (p_0[0]), .B (p_1[0]));
INV_X1 slo__sro_c5 (.ZN (slo__sro_n71), .A (n_29));
NAND2_X1 slo__sro_c6 (.ZN (slo__sro_n70), .A1 (p_0[29]), .A2 (p_1[29]));
NOR2_X1 slo__sro_c7 (.ZN (slo__sro_n69), .A1 (p_1[29]), .A2 (p_0[29]));
OAI21_X2 slo__sro_c8 (.ZN (slo__sro_n68), .A (slo__sro_n70), .B1 (slo__sro_n71), .B2 (slo__sro_n69));
XNOR2_X1 slo__sro_c9 (.ZN (slo__sro_n67), .A (p_1[29]), .B (p_0[29]));
XNOR2_X1 slo__sro_c10 (.ZN (p_2[29]), .A (n_29), .B (slo__sro_n67));
NAND2_X1 slo__sro_c46 (.ZN (slo__sro_n110), .A1 (p_1[17]), .A2 (p_0[17]));
NOR2_X1 slo__sro_c47 (.ZN (slo__sro_n109), .A1 (p_1[17]), .A2 (p_0[17]));
OAI21_X1 slo__sro_c48 (.ZN (n_18), .A (slo__sro_n110), .B1 (slo__sro_n111), .B2 (slo__sro_n109));
XNOR2_X1 slo__sro_c49 (.ZN (slo__sro_n108), .A (p_1[17]), .B (p_0[17]));
XNOR2_X1 slo__sro_c50 (.ZN (p_2[17]), .A (slo__sro_n108), .B (n_17));
NAND2_X1 slo__sro_c60 (.ZN (slo__sro_n123), .A1 (p_1[15]), .A2 (p_0[15]));
NOR2_X1 slo__sro_c61 (.ZN (slo__sro_n122), .A1 (p_1[15]), .A2 (p_0[15]));
OAI21_X2 slo__sro_c62 (.ZN (n_16), .A (slo__sro_n123), .B1 (slo__sro_n124), .B2 (slo__sro_n122));
XNOR2_X1 slo__sro_c63 (.ZN (slo__sro_n121), .A (p_1[15]), .B (p_0[15]));
XNOR2_X1 slo__sro_c64 (.ZN (p_2[15]), .A (slo__sro_n195), .B (slo__sro_n121));
NAND2_X1 slo__sro_c87 (.ZN (slo__sro_n151), .A1 (p_1[7]), .A2 (p_0[7]));
NOR2_X1 slo__sro_c88 (.ZN (slo__sro_n150), .A1 (p_1[7]), .A2 (p_0[7]));
OAI21_X1 slo__sro_c89 (.ZN (n_8), .A (slo__sro_n151), .B1 (slo__sro_n152), .B2 (slo__sro_n150));
XNOR2_X1 slo__sro_c90 (.ZN (slo__sro_n149), .A (p_1[7]), .B (p_0[7]));
XNOR2_X1 slo__sro_c91 (.ZN (p_2[7]), .A (slo__sro_n149), .B (n_7));
NAND2_X1 slo__sro_c114 (.ZN (slo__sro_n179), .A1 (n_24), .A2 (p_0[24]));
NAND2_X1 slo__sro_c115 (.ZN (slo__sro_n178), .A1 (n_24), .A2 (p_1[24]));
NAND3_X1 slo__sro_c116 (.ZN (n_25), .A1 (slo__sro_n180), .A2 (slo__sro_n178), .A3 (slo__sro_n179));
XNOR2_X1 slo__sro_c117 (.ZN (slo__sro_n177), .A (p_1[24]), .B (p_0[24]));
XNOR2_X1 slo__sro_c118 (.ZN (p_2[24]), .A (slo__sro_n177), .B (n_24));
NAND2_X1 slo__sro_c132 (.ZN (slo__sro_n197), .A1 (p_1[14]), .A2 (p_0[14]));
NOR2_X1 slo__sro_c133 (.ZN (slo__sro_n196), .A1 (p_1[14]), .A2 (p_0[14]));
OAI21_X2 slo__sro_c134 (.ZN (slo__sro_n195), .A (slo__sro_n197), .B1 (slo__sro_n198), .B2 (slo__sro_n196));
XNOR2_X1 slo__sro_c135 (.ZN (slo__sro_n194), .A (p_1[14]), .B (p_0[14]));
XNOR2_X1 slo__sro_c136 (.ZN (p_2[14]), .A (n_14), .B (slo__sro_n194));
NAND2_X1 slo__sro_c208 (.ZN (slo__sro_n269), .A1 (p_1[10]), .A2 (p_0[10]));
NOR2_X2 slo__sro_c209 (.ZN (slo__sro_n268), .A1 (p_1[10]), .A2 (p_0[10]));
OAI21_X1 slo__sro_c210 (.ZN (slo__sro_n267), .A (slo__sro_n269), .B1 (slo__sro_n270), .B2 (slo__sro_n268));
XNOR2_X1 slo__sro_c211 (.ZN (slo__sro_n266), .A (p_1[10]), .B (p_0[10]));
XNOR2_X1 slo__sro_c212 (.ZN (p_2[10]), .A (slo__sro_n266), .B (n_10));
NAND2_X1 slo__sro_c222 (.ZN (slo__sro_n286), .A1 (p_1[22]), .A2 (p_0[22]));
NOR2_X1 slo__sro_c223 (.ZN (slo__sro_n285), .A1 (p_1[22]), .A2 (p_0[22]));
OAI21_X2 slo__sro_c224 (.ZN (slo__sro_n284), .A (slo__sro_n286), .B1 (slo__sro_n287), .B2 (slo__sro_n285));
XNOR2_X1 slo__sro_c225 (.ZN (slo__sro_n283), .A (p_1[22]), .B (p_0[22]));
XNOR2_X1 slo__sro_c226 (.ZN (p_2[22]), .A (slo__sro_n283), .B (n_22));
NOR2_X1 slo__sro_c244 (.ZN (slo__sro_n314), .A1 (n_33), .A2 (p_0[30]));
NAND2_X1 slo__sro_c245 (.ZN (slo__sro_n313), .A1 (slo__sro_n315), .A2 (slo__sro_n314));
NOR2_X1 slo__sro_c246 (.ZN (slo__sro_n312), .A1 (p_1[30]), .A2 (n_34));
INV_X1 slo__sro_c247 (.ZN (slo__sro_n311), .A (slo__sro_n312));
OAI21_X2 slo__sro_c248 (.ZN (slo__sro_n310), .A (slo__sro_n313), .B1 (n_32), .B2 (slo__sro_n311));
INV_X1 slo__sro_c414 (.ZN (slo__sro_n551), .A (n_16));
INV_X1 slo__sro_c333 (.ZN (slo__sro_n456), .A (n_28));
NOR2_X1 slo__sro_c335 (.ZN (slo__sro_n454), .A1 (p_1[28]), .A2 (p_0[28]));
INV_X1 slo__sro_c315 (.ZN (slo__sro_n436), .A (n_20));
NAND2_X1 slo__sro_c316 (.ZN (slo__sro_n435), .A1 (p_1[20]), .A2 (p_0[20]));
NOR2_X1 slo__sro_c317 (.ZN (slo__sro_n434), .A1 (p_1[20]), .A2 (p_0[20]));
OAI21_X1 slo__sro_c318 (.ZN (slo__sro_n433), .A (slo__sro_n435), .B1 (slo__sro_n436), .B2 (slo__sro_n434));
XNOR2_X1 slo__sro_c319 (.ZN (slo__sro_n432), .A (p_1[20]), .B (p_0[20]));
XNOR2_X1 slo__sro_c320 (.ZN (p_2[20]), .A (slo__sro_n432), .B (n_20));
XNOR2_X2 slo__sro_c337 (.ZN (slo__sro_n453), .A (p_1[28]), .B (p_0[28]));
XNOR2_X1 slo__sro_c338 (.ZN (p_2[28]), .A (n_28), .B (slo__sro_n453));
NOR2_X1 slo__sro_c416 (.ZN (slo__sro_n549), .A1 (p_1[16]), .A2 (p_0[16]));
OAI21_X1 slo__sro_c417 (.ZN (n_17), .A (slo__sro_n550), .B1 (slo__sro_n551), .B2 (slo__sro_n549));
XNOR2_X1 slo__sro_c418 (.ZN (slo__sro_n548), .A (p_1[16]), .B (p_0[16]));
XNOR2_X1 slo__sro_c419 (.ZN (p_2[16]), .A (n_16), .B (slo__sro_n548));
OAI21_X1 CLOCK_slo__c1187 (.ZN (CLOCK_slo__n1670), .A (slo__sro_n550), .B1 (slo__sro_n551), .B2 (slo__sro_n549));
OAI21_X2 CLOCK_slo__sro_c927 (.ZN (n_10), .A (CLOCK_slo__sro_n1431), .B1 (CLOCK_slo__sro_n1432), .B2 (CLOCK_slo__sro_n1430));
XNOR2_X1 CLOCK_slo__sro_c928 (.ZN (CLOCK_slo__sro_n1429), .A (p_1[9]), .B (p_0[9]));
INV_X1 slo__sro_c538 (.ZN (slo__sro_n754), .A (n_19));
NAND2_X1 slo__sro_c539 (.ZN (slo__sro_n753), .A1 (p_1[19]), .A2 (p_0[19]));
NOR2_X1 slo__sro_c540 (.ZN (slo__sro_n752), .A1 (p_1[19]), .A2 (p_0[19]));
OAI21_X1 slo__sro_c541 (.ZN (n_20), .A (slo__sro_n753), .B1 (slo__sro_n754), .B2 (slo__sro_n752));
XNOR2_X1 slo__sro_c542 (.ZN (slo__sro_n751), .A (p_1[19]), .B (p_0[19]));
XNOR2_X1 slo__sro_c543 (.ZN (p_2[19]), .A (n_19), .B (slo__sro_n751));
INV_X1 CLOCK_slo__sro_c924 (.ZN (CLOCK_slo__sro_n1432), .A (n_9));
NAND2_X1 CLOCK_slo__sro_c925 (.ZN (CLOCK_slo__sro_n1431), .A1 (p_1[9]), .A2 (p_0[9]));
NOR2_X2 CLOCK_slo__sro_c926 (.ZN (CLOCK_slo__sro_n1430), .A1 (p_1[9]), .A2 (p_0[9]));
INV_X1 CLOCK_slo__sro_c984 (.ZN (CLOCK_slo__sro_n1486), .A (p_1[8]));
INV_X1 CLOCK_slo__sro_c951 (.ZN (CLOCK_slo__sro_n1457), .A (n_27));
NAND2_X1 CLOCK_slo__sro_c952 (.ZN (CLOCK_slo__sro_n1456), .A1 (p_1[27]), .A2 (p_0[27]));
NOR2_X1 CLOCK_slo__sro_c953 (.ZN (CLOCK_slo__sro_n1455), .A1 (p_1[27]), .A2 (p_0[27]));
OAI21_X2 CLOCK_slo__sro_c954 (.ZN (n_28), .A (CLOCK_slo__sro_n1456), .B1 (CLOCK_slo__sro_n1457), .B2 (CLOCK_slo__sro_n1455));
XNOR2_X1 CLOCK_slo__sro_c955 (.ZN (CLOCK_slo__sro_n1454), .A (p_1[27]), .B (p_0[27]));
XNOR2_X1 CLOCK_slo__sro_c956 (.ZN (p_2[27]), .A (CLOCK_slo__sro_n1454), .B (n_27));
NAND2_X1 CLOCK_slo__sro_c986 (.ZN (CLOCK_slo__sro_n1484), .A1 (CLOCK_slo__sro_n1487), .A2 (CLOCK_slo__sro_n1486));
NAND2_X1 CLOCK_slo__sro_c987 (.ZN (CLOCK_slo__sro_n1483), .A1 (n_8), .A2 (CLOCK_slo__sro_n1484));
NAND2_X1 CLOCK_slo__sro_c988 (.ZN (n_9), .A1 (CLOCK_slo__sro_n1483), .A2 (CLOCK_slo__sro_n1485));
XNOR2_X1 CLOCK_slo__sro_c989 (.ZN (CLOCK_slo__sro_n1482), .A (p_1[8]), .B (p_0[8]));
XNOR2_X1 CLOCK_slo__sro_c990 (.ZN (p_2[8]), .A (n_8), .B (CLOCK_slo__sro_n1482));
NAND2_X1 CLOCK_slo__sro_c1127 (.ZN (CLOCK_slo__sro_n1625), .A1 (p_0[23]), .A2 (p_1[23]));
OAI21_X1 CLOCK_slo__sro_c1128 (.ZN (CLOCK_slo__sro_n1624), .A (slo__sro_n284), .B1 (p_1[23]), .B2 (p_0[23]));
NAND2_X1 CLOCK_slo__sro_c1129 (.ZN (n_24), .A1 (CLOCK_slo__sro_n1624), .A2 (CLOCK_slo__sro_n1625));
XNOR2_X1 CLOCK_slo__sro_c1130 (.ZN (CLOCK_slo__sro_n1623), .A (p_1[23]), .B (p_0[23]));
XNOR2_X1 CLOCK_slo__sro_c1131 (.ZN (p_2[23]), .A (CLOCK_slo__sro_n1623), .B (slo__sro_n284));

endmodule //datapath__0_237

module datapath__0_236 (p_0_25_PP_0, Multiplier, p_0, p_1);

output [31:0] p_1;
input [31:0] Multiplier;
input [31:0] p_0;
input p_0_25_PP_0;
wire slo_n354;
wire CLOCK_slo__sro_n1651;
wire slo__sro_n626;
wire n_1;
wire n_2;
wire n_3;
wire n_4;
wire n_5;
wire n_6;
wire n_8;
wire n_9;
wire n_11;
wire n_12;
wire n_16;
wire n_17;
wire CLOCK_slo__sro_n1648;
wire n_19;
wire n_20;
wire n_22;
wire n_25;
wire n_27;
wire n_30;
wire n_32;
wire n_34;
wire n_33;
wire slo__sro_n1115;
wire slo__sro_n59;
wire slo__sro_n60;
wire slo__sro_n61;
wire slo__sro_n72;
wire slo__sro_n73;
wire slo__sro_n74;
wire slo__sro_n75;
wire slo__sro_n76;
wire slo__sro_n91;
wire slo__sro_n92;
wire slo__sro_n93;
wire slo__sro_n94;
wire slo__sro_n106;
wire slo__sro_n107;
wire slo__sro_n108;
wire slo__n846;
wire slo__sro_n150;
wire slo__sro_n151;
wire slo__sro_n152;
wire slo__sro_n132;
wire slo__sro_n133;
wire slo__sro_n134;
wire slo__sro_n135;
wire slo__sro_n136;
wire slo__sro_n162;
wire slo__sro_n163;
wire slo__sro_n164;
wire slo__sro_n165;
wire slo__sro_n175;
wire slo__sro_n176;
wire slo__sro_n177;
wire slo__sro_n178;
wire slo__sro_n196;
wire slo__sro_n197;
wire slo__sro_n198;
wire slo__sro_n199;
wire slo__sro_n200;
wire slo__sro_n213;
wire slo__sro_n214;
wire slo__sro_n215;
wire slo__sro_n216;
wire slo__sro_n228;
wire slo__sro_n229;
wire slo__sro_n230;
wire slo__sro_n243;
wire slo__sro_n244;
wire slo__sro_n245;
wire slo__sro_n246;
wire slo__sro_n247;
wire slo__sro_n262;
wire slo__sro_n263;
wire slo__sro_n264;
wire slo__sro_n265;
wire slo__sro_n266;
wire slo__sro_n267;
wire slo__sro_n268;
wire slo__sro_n283;
wire slo__sro_n284;
wire slo__sro_n285;
wire slo__sro_n286;
wire slo___n336;
wire slo__n315;
wire slo__sro_n623;
wire slo__n482;
wire slo__sro_n624;
wire slo__sro_n625;
wire slo__sro_n450;
wire slo__sro_n451;
wire slo__sro_n452;
wire slo__sro_n453;
wire slo__sro_n627;
wire slo__mro_n776;
wire slo__sro_n858;
wire slo__n533;
wire slo__sro_n859;
wire slo__sro_n860;
wire slo__sro_n861;
wire slo__sro_n922;
wire slo__sro_n923;
wire slo__sro_n924;
wire slo__sro_n925;
wire slo__sro_n926;
wire slo__sro_n966;
wire slo__sro_n967;
wire slo__sro_n968;
wire slo__sro_n969;
wire slo__sro_n970;
wire slo__mro_n1026;
wire slo__mro_n1027;
wire slo__mro_n1028;
wire slo__mro_n1029;
wire slo__mro_n1030;
wire CLOCK_slo__sro_n1650;
wire CLOCK_slo__sro_n2040;
wire CLOCK_slo__sro_n1647;
wire CLOCK_slo__sro_n1649;
wire CLOCK_slo__sro_n1652;
wire CLOCK_slo__mro_n1687;


INV_X1 i_36 (.ZN (n_34), .A (Multiplier[30]));
INV_X1 i_35 (.ZN (n_33), .A (p_0[30]));
INV_X2 i_34 (.ZN (n_32), .A (n_30));
OAI22_X1 CLOCK_slo__sro_c1587 (.ZN (CLOCK_slo__sro_n2040), .A1 (n_33), .A2 (Multiplier[30])
    , .B1 (p_0[30]), .B2 (n_34));
XNOR2_X1 i_0 (.ZN (p_1[30]), .A (CLOCK_slo__sro_n2040), .B (n_32));
NAND2_X1 slo__sro_c49 (.ZN (slo__sro_n108), .A1 (slo__sro_n73), .A2 (Multiplier[7]));
INV_X1 slo__sro_c193 (.ZN (slo__sro_n268), .A (Multiplier[27]));
INV_X1 slo__sro_c211 (.ZN (slo__sro_n286), .A (slo__sro_n624));
INV_X2 slo__sro_c177 (.ZN (slo__sro_n247), .A (slo__sro_n263));
INV_X1 slo__sro_c137 (.ZN (slo__sro_n200), .A (slo__n482));
INV_X1 slo__sro_c102 (.ZN (slo__sro_n165), .A (slo__sro_n450));
INV_X1 slo__sro_c689 (.ZN (slo__sro_n970), .A (n_9));
NAND2_X2 slo__sro_c163 (.ZN (slo__sro_n230), .A1 (slo__sro_n176), .A2 (Multiplier[26]));
NAND2_X1 slo__sro_c116 (.ZN (slo__sro_n178), .A1 (n_25), .A2 (Multiplier[25]));
OAI21_X2 slo__sro_c455 (.ZN (slo__sro_n624), .A (slo__sro_n626), .B1 (slo__sro_n627), .B2 (slo__sro_n625));
FA_X1 i_20 (.CO (n_20), .S (p_1[19]), .A (Multiplier[19]), .B (p_0[19]), .CI (n_19));
FA_X1 i_19 (.CO (n_19), .S (p_1[18]), .A (Multiplier[18]), .B (p_0[18]), .CI (slo__sro_n1115));
INV_X2 slo__sro_c17 (.ZN (slo__sro_n76), .A (n_6));
INV_X1 CLOCK_slo__mro_c1174 (.ZN (slo__mro_n1030), .A (n_32));
INV_X1 slo___L2_c2_c248 (.ZN (slo_n354), .A (p_0[25]));
XNOR2_X2 slo__mro_c531 (.ZN (slo__mro_n776), .A (slo__sro_n923), .B (Multiplier[24]));
NAND2_X1 slo__sro_c151 (.ZN (slo__sro_n216), .A1 (n_22), .A2 (Multiplier[22]));
NAND2_X1 slo__sro_c103 (.ZN (slo__sro_n164), .A1 (p_0[21]), .A2 (Multiplier[21]));
INV_X2 slo__sro_c654 (.ZN (slo__sro_n926), .A (slo__sro_n214));
FA_X1 i_11 (.CO (n_11), .S (p_1[10]), .A (Multiplier[10]), .B (p_0[10]), .CI (slo__sro_n967));
XNOR2_X1 CLOCK_slo__mro_c1186 (.ZN (CLOCK_slo__mro_n1687), .A (p_0[20]), .B (Multiplier[20]));
FA_X1 i_9 (.CO (n_9), .S (p_1[8]), .A (Multiplier[8]), .B (p_0[8]), .CI (n_8));
INV_X1 slo__sro_c88 (.ZN (slo__sro_n152), .A (slo__sro_n923));
INV_X2 slo__sro_c33 (.ZN (slo__sro_n94), .A (slo__sro_n244));
FA_X1 i_6 (.CO (n_6), .S (p_1[5]), .A (Multiplier[5]), .B (p_0[5]), .CI (n_5));
FA_X1 i_5 (.CO (n_5), .S (p_1[4]), .A (Multiplier[4]), .B (p_0[4]), .CI (n_4));
FA_X1 i_4 (.CO (n_4), .S (p_1[3]), .A (Multiplier[3]), .B (p_0[3]), .CI (n_3));
FA_X1 i_3 (.CO (n_3), .S (p_1[2]), .A (Multiplier[2]), .B (p_0[2]), .CI (n_2));
FA_X1 i_2 (.CO (n_2), .S (p_1[1]), .A (Multiplier[1]), .B (p_0[1]), .CI (n_1));
HA_X1 i_1 (.CO (n_1), .S (p_1[0]), .A (Multiplier[0]), .B (p_0[0]));
INV_X1 slo__sro_c605 (.ZN (slo__sro_n861), .A (n_11));
NAND2_X1 slo__sro_c4 (.ZN (slo__sro_n61), .A1 (p_0[17]), .A2 (Multiplier[17]));
NOR2_X2 slo__sro_c5 (.ZN (slo__sro_n60), .A1 (p_0[17]), .A2 (Multiplier[17]));
NAND2_X1 CLOCK_slo__sro_c1139 (.ZN (CLOCK_slo__sro_n1649), .A1 (CLOCK_slo__sro_n1652), .A2 (CLOCK_slo__sro_n1651));
XNOR2_X1 slo__sro_c7 (.ZN (slo__sro_n59), .A (p_0[17]), .B (Multiplier[17]));
XNOR2_X1 slo__sro_c8 (.ZN (p_1[17]), .A (slo__sro_n59), .B (n_17));
NAND2_X1 slo__sro_c18 (.ZN (slo__sro_n75), .A1 (p_0[6]), .A2 (Multiplier[6]));
NOR2_X2 slo__sro_c19 (.ZN (slo__sro_n74), .A1 (p_0[6]), .A2 (Multiplier[6]));
OAI21_X2 slo__sro_c20 (.ZN (slo__sro_n73), .A (slo__sro_n75), .B1 (slo__sro_n76), .B2 (slo__sro_n74));
XNOR2_X1 slo__sro_c21 (.ZN (slo__sro_n72), .A (p_0[6]), .B (Multiplier[6]));
XNOR2_X1 slo__sro_c22 (.ZN (p_1[6]), .A (slo__sro_n72), .B (n_6));
NAND2_X1 slo__sro_c34 (.ZN (slo__sro_n93), .A1 (p_0[29]), .A2 (Multiplier[29]));
NOR2_X1 slo__sro_c35 (.ZN (slo__sro_n92), .A1 (p_0[29]), .A2 (Multiplier[29]));
OAI21_X2 slo__sro_c36 (.ZN (n_30), .A (slo__sro_n93), .B1 (slo__sro_n92), .B2 (slo__sro_n94));
XNOR2_X2 slo__sro_c37 (.ZN (slo__sro_n91), .A (p_0[29]), .B (Multiplier[29]));
XNOR2_X2 slo__sro_c38 (.ZN (p_1[29]), .A (slo__sro_n91), .B (slo__sro_n244));
OAI21_X1 slo__sro_c50 (.ZN (slo__sro_n107), .A (p_0[7]), .B1 (slo__sro_n73), .B2 (Multiplier[7]));
NAND2_X1 slo__sro_c51 (.ZN (n_8), .A1 (slo__sro_n107), .A2 (slo__sro_n108));
XNOR2_X2 slo__sro_c52 (.ZN (slo__sro_n106), .A (slo__n315), .B (Multiplier[7]));
XNOR2_X2 slo__sro_c53 (.ZN (p_1[7]), .A (slo__sro_n106), .B (p_0[7]));
NAND2_X1 slo__sro_c89 (.ZN (slo__sro_n151), .A1 (p_0[24]), .A2 (Multiplier[24]));
NOR2_X2 slo__sro_c90 (.ZN (slo__sro_n150), .A1 (p_0[24]), .A2 (Multiplier[24]));
OAI21_X2 slo__sro_c91 (.ZN (n_25), .A (slo__sro_n151), .B1 (slo__sro_n150), .B2 (slo__sro_n152));
INV_X1 slo__L1_c595 (.ZN (slo__n846), .A (n_17));
INV_X1 slo__sro_c74 (.ZN (slo__sro_n136), .A (n_12));
NAND2_X1 slo__sro_c75 (.ZN (slo__sro_n135), .A1 (p_0[12]), .A2 (Multiplier[12]));
NOR2_X1 slo__sro_c76 (.ZN (slo__sro_n134), .A1 (p_0[12]), .A2 (Multiplier[12]));
OAI21_X1 slo__sro_c77 (.ZN (slo__sro_n133), .A (slo__sro_n135), .B1 (slo__sro_n136), .B2 (slo__sro_n134));
XNOR2_X2 slo__sro_c78 (.ZN (slo__sro_n132), .A (p_0[12]), .B (Multiplier[12]));
XNOR2_X2 slo__sro_c79 (.ZN (p_1[12]), .A (slo__sro_n132), .B (n_12));
NOR2_X2 slo__sro_c104 (.ZN (slo__sro_n163), .A1 (p_0[21]), .A2 (Multiplier[21]));
OAI21_X2 slo__sro_c105 (.ZN (n_22), .A (slo__sro_n164), .B1 (slo__sro_n163), .B2 (slo__sro_n165));
XNOR2_X1 slo__sro_c106 (.ZN (slo__sro_n162), .A (p_0[21]), .B (Multiplier[21]));
XNOR2_X1 slo__sro_c107 (.ZN (p_1[21]), .A (slo__sro_n162), .B (slo__sro_n450));
OAI21_X2 slo__sro_c117 (.ZN (slo__sro_n177), .A (slo_n354), .B1 (n_25), .B2 (Multiplier[25]));
NAND2_X4 slo__sro_c118 (.ZN (slo__sro_n176), .A1 (slo__sro_n177), .A2 (slo__sro_n178));
XNOR2_X1 slo__sro_c119 (.ZN (slo__sro_n175), .A (n_25), .B (Multiplier[25]));
XNOR2_X1 slo__sro_c120 (.ZN (p_1[25]), .A (slo__sro_n175), .B (slo___n336));
NAND2_X1 slo__sro_c138 (.ZN (slo__sro_n199), .A1 (p_0[13]), .A2 (Multiplier[13]));
NOR2_X2 slo__sro_c139 (.ZN (slo__sro_n198), .A1 (p_0[13]), .A2 (Multiplier[13]));
OAI21_X2 slo__sro_c140 (.ZN (slo__sro_n197), .A (slo__sro_n199), .B1 (slo__sro_n200), .B2 (slo__sro_n198));
XNOR2_X1 slo__sro_c141 (.ZN (slo__sro_n196), .A (p_0[13]), .B (Multiplier[13]));
XNOR2_X1 slo__sro_c142 (.ZN (p_1[13]), .A (slo__sro_n196), .B (slo__sro_n133));
OAI21_X1 slo__sro_c152 (.ZN (slo__sro_n215), .A (p_0[22]), .B1 (n_22), .B2 (Multiplier[22]));
NAND2_X2 slo__sro_c153 (.ZN (slo__sro_n214), .A1 (slo__sro_n215), .A2 (slo__sro_n216));
XNOR2_X2 slo__sro_c154 (.ZN (slo__sro_n213), .A (n_22), .B (Multiplier[22]));
XNOR2_X2 slo__sro_c155 (.ZN (p_1[22]), .A (slo__sro_n213), .B (p_0[22]));
OAI21_X2 slo__sro_c164 (.ZN (slo__sro_n229), .A (p_0[26]), .B1 (slo__sro_n176), .B2 (Multiplier[26]));
NAND2_X2 slo__sro_c165 (.ZN (n_27), .A1 (slo__sro_n229), .A2 (slo__sro_n230));
XNOR2_X1 slo__sro_c166 (.ZN (slo__sro_n228), .A (slo__sro_n176), .B (Multiplier[26]));
XNOR2_X1 slo__sro_c167 (.ZN (p_1[26]), .A (slo__sro_n228), .B (p_0[26]));
NAND2_X1 slo__sro_c178 (.ZN (slo__sro_n246), .A1 (p_0[28]), .A2 (Multiplier[28]));
NOR2_X2 slo__sro_c179 (.ZN (slo__sro_n245), .A1 (p_0[28]), .A2 (Multiplier[28]));
OAI21_X4 slo__sro_c180 (.ZN (slo__sro_n244), .A (slo__sro_n246), .B1 (slo__sro_n247), .B2 (slo__sro_n245));
XNOR2_X2 slo__sro_c181 (.ZN (slo__sro_n243), .A (p_0[28]), .B (Multiplier[28]));
XNOR2_X1 slo__sro_c182 (.ZN (p_1[28]), .A (slo__sro_n243), .B (slo__sro_n263));
INV_X1 slo__sro_c194 (.ZN (slo__sro_n267), .A (n_27));
NAND2_X1 slo__sro_c195 (.ZN (slo__sro_n266), .A1 (n_27), .A2 (Multiplier[27]));
NAND2_X1 slo__sro_c196 (.ZN (slo__sro_n265), .A1 (slo__sro_n267), .A2 (slo__sro_n268));
NAND2_X1 slo__sro_c197 (.ZN (slo__sro_n264), .A1 (slo__sro_n265), .A2 (p_0[27]));
NAND2_X1 slo__sro_c198 (.ZN (slo__sro_n263), .A1 (slo__sro_n264), .A2 (slo__sro_n266));
XNOR2_X2 slo__sro_c199 (.ZN (slo__sro_n262), .A (slo__n533), .B (Multiplier[27]));
XNOR2_X1 slo__sro_c200 (.ZN (p_1[27]), .A (slo__sro_n262), .B (p_0[27]));
NAND2_X1 slo__sro_c212 (.ZN (slo__sro_n285), .A1 (p_0[15]), .A2 (Multiplier[15]));
NOR2_X2 slo__sro_c213 (.ZN (slo__sro_n284), .A1 (p_0[15]), .A2 (Multiplier[15]));
OAI21_X1 slo__sro_c214 (.ZN (n_16), .A (slo__sro_n285), .B1 (slo__sro_n284), .B2 (slo__sro_n286));
XNOR2_X1 slo__sro_c215 (.ZN (slo__sro_n283), .A (p_0[15]), .B (Multiplier[15]));
XNOR2_X1 slo__sro_c216 (.ZN (p_1[15]), .A (slo__sro_n283), .B (slo__sro_n624));
INV_X1 slo___L2_c3_c249 (.ZN (slo___n336), .A (p_0_25_PP_0));
NAND2_X1 slo__sro_c453 (.ZN (slo__sro_n626), .A1 (p_0[14]), .A2 (Multiplier[14]));
OAI21_X2 slo__c237 (.ZN (slo__n315), .A (slo__sro_n75), .B1 (slo__sro_n76), .B2 (slo__sro_n74));
INV_X1 slo__sro_c452 (.ZN (slo__sro_n627), .A (slo__sro_n197));
OAI21_X1 slo__c330 (.ZN (slo__n482), .A (slo__sro_n135), .B1 (slo__sro_n134), .B2 (slo__sro_n136));
NOR2_X2 slo__sro_c454 (.ZN (slo__sro_n625), .A1 (p_0[14]), .A2 (Multiplier[14]));
INV_X2 slo__sro_c305 (.ZN (slo__sro_n453), .A (n_20));
NAND2_X1 slo__sro_c306 (.ZN (slo__sro_n452), .A1 (p_0[20]), .A2 (Multiplier[20]));
NOR2_X1 slo__sro_c307 (.ZN (slo__sro_n451), .A1 (p_0[20]), .A2 (Multiplier[20]));
OAI21_X2 slo__sro_c308 (.ZN (slo__sro_n450), .A (slo__sro_n452), .B1 (slo__sro_n453), .B2 (slo__sro_n451));
OAI21_X1 CLOCK_slo__sro_c1311 (.ZN (slo__sro_n1115), .A (slo__sro_n61), .B1 (slo__sro_n60), .B2 (slo__n846));
XNOR2_X1 slo__sro_c456 (.ZN (slo__sro_n623), .A (p_0[14]), .B (Multiplier[14]));
XNOR2_X1 slo__sro_c457 (.ZN (p_1[14]), .A (slo__sro_n623), .B (slo__sro_n197));
XNOR2_X2 slo__mro_c532 (.ZN (p_1[24]), .A (slo__mro_n776), .B (p_0[24]));
NAND2_X1 slo__sro_c606 (.ZN (slo__sro_n860), .A1 (p_0[11]), .A2 (Multiplier[11]));
NOR2_X1 slo__sro_c607 (.ZN (slo__sro_n859), .A1 (p_0[11]), .A2 (Multiplier[11]));
NAND2_X2 slo__c370 (.ZN (slo__n533), .A1 (slo__sro_n229), .A2 (slo__sro_n230));
OAI21_X2 slo__sro_c608 (.ZN (n_12), .A (slo__sro_n860), .B1 (slo__sro_n861), .B2 (slo__sro_n859));
XNOR2_X1 slo__sro_c609 (.ZN (slo__sro_n858), .A (p_0[11]), .B (Multiplier[11]));
XNOR2_X1 slo__sro_c610 (.ZN (p_1[11]), .A (slo__sro_n858), .B (n_11));
NAND2_X1 slo__sro_c655 (.ZN (slo__sro_n925), .A1 (p_0[23]), .A2 (Multiplier[23]));
NOR2_X1 slo__sro_c656 (.ZN (slo__sro_n924), .A1 (p_0[23]), .A2 (Multiplier[23]));
OAI21_X2 slo__sro_c657 (.ZN (slo__sro_n923), .A (slo__sro_n925), .B1 (slo__sro_n926), .B2 (slo__sro_n924));
XNOR2_X2 slo__sro_c658 (.ZN (slo__sro_n922), .A (p_0[23]), .B (Multiplier[23]));
XNOR2_X2 slo__sro_c659 (.ZN (p_1[23]), .A (slo__sro_n922), .B (slo__sro_n214));
NAND2_X1 slo__sro_c690 (.ZN (slo__sro_n969), .A1 (p_0[9]), .A2 (Multiplier[9]));
NOR2_X1 slo__sro_c691 (.ZN (slo__sro_n968), .A1 (p_0[9]), .A2 (Multiplier[9]));
OAI21_X2 slo__sro_c692 (.ZN (slo__sro_n967), .A (slo__sro_n969), .B1 (slo__sro_n970), .B2 (slo__sro_n968));
XNOR2_X1 slo__sro_c693 (.ZN (slo__sro_n966), .A (p_0[9]), .B (Multiplier[9]));
XNOR2_X1 slo__sro_c694 (.ZN (p_1[9]), .A (slo__sro_n966), .B (n_9));
INV_X1 slo__mro_c736 (.ZN (slo__mro_n1029), .A (Multiplier[30]));
NOR2_X1 slo__mro_c737 (.ZN (slo__mro_n1028), .A1 (n_30), .A2 (n_33));
NOR2_X1 slo__mro_c738 (.ZN (slo__mro_n1027), .A1 (p_0[30]), .A2 (n_34));
XNOR2_X1 CLOCK_slo__mro_c1187 (.ZN (p_1[20]), .A (CLOCK_slo__mro_n1687), .B (n_20));
XNOR2_X1 CLOCK_slo__sro_c1143 (.ZN (p_1[16]), .A (n_16), .B (CLOCK_slo__sro_n1647));
XNOR2_X1 CLOCK_slo__sro_c1142 (.ZN (CLOCK_slo__sro_n1647), .A (p_0[16]), .B (Multiplier[16]));
NAND2_X1 CLOCK_slo__sro_c1138 (.ZN (CLOCK_slo__sro_n1650), .A1 (p_0[16]), .A2 (Multiplier[16]));
INV_X1 CLOCK_slo__sro_c1136 (.ZN (CLOCK_slo__sro_n1652), .A (Multiplier[16]));
INV_X1 CLOCK_slo__sro_c1137 (.ZN (CLOCK_slo__sro_n1651), .A (p_0[16]));
NAND2_X1 CLOCK_slo__sro_c1140 (.ZN (CLOCK_slo__sro_n1648), .A1 (CLOCK_slo__sro_n1649), .A2 (n_16));
NAND2_X2 CLOCK_slo__sro_c1141 (.ZN (n_17), .A1 (CLOCK_slo__sro_n1648), .A2 (CLOCK_slo__sro_n1650));
AOI22_X2 CLOCK_slo__mro_c1175 (.ZN (slo__mro_n1026), .A1 (slo__mro_n1030), .A2 (slo__mro_n1027)
    , .B1 (slo__mro_n1028), .B2 (slo__mro_n1029));
XNOR2_X2 CLOCK_slo__mro_c1176 (.ZN (p_1[31]), .A (slo__mro_n1026), .B (Multiplier[31]));

endmodule //datapath__0_236

module datapath__0_232 (p_0, p_1, p_2);

output [31:0] p_2;
input [31:0] p_0;
input [31:0] p_1;
wire spw_n2396;
wire slo__sro_n594;
wire n_1;
wire n_2;
wire n_3;
wire n_5;
wire CLOCK_slo__sro_n1762;
wire n_7;
wire n_8;
wire n_9;
wire n_10;
wire slo__sro_n390;
wire n_12;
wire n_14;
wire CLOCK_slo__sro_n1635;
wire n_17;
wire slo__sro_n841;
wire slo__sro_n1028;
wire slo__sro_n589;
wire n_21;
wire n_22;
wire n_24;
wire n_25;
wire n_26;
wire n_27;
wire n_28;
wire n_29;
wire n_30;
wire n_32;
wire n_0;
wire n_34;
wire n_33;
wire n_31;
wire slo__sro_n253;
wire slo__sro_n254;
wire slo__sro_n255;
wire slo__sro_n256;
wire slo__sro_n73;
wire slo__sro_n74;
wire slo__sro_n75;
wire slo__sro_n76;
wire slo__sro_n101;
wire slo__sro_n102;
wire slo__sro_n103;
wire slo__sro_n104;
wire slo__sro_n127;
wire slo__sro_n128;
wire slo__sro_n129;
wire CLOCK_slo__sro_n1636;
wire slo__sro_n270;
wire slo__sro_n271;
wire slo__sro_n272;
wire slo__sro_n273;
wire slo__sro_n274;
wire slo__sro_n590;
wire slo__sro_n591;
wire slo__sro_n592;
wire slo__sro_n593;
wire slo__sro_n301;
wire slo__sro_n302;
wire slo__sro_n303;
wire slo__sro_n304;
wire slo__sro_n305;
wire slo__sro_n388;
wire slo__sro_n389;
wire slo__sro_n343;
wire slo__sro_n344;
wire slo__sro_n345;
wire slo__sro_n346;
wire slo__sro_n347;
wire slo__sro_n391;
wire slo__sro_n838;
wire slo__sro_n839;
wire slo__sro_n840;
wire slo__sro_n720;
wire slo__sro_n721;
wire slo__sro_n723;
wire slo__sro_n1029;
wire slo__sro_n1014;
wire slo__sro_n1015;
wire slo__sro_n1016;
wire slo__sro_n1017;
wire slo__sro_n1026;
wire slo__sro_n1027;
wire CLOCK_slo__sro_n1637;
wire CLOCK_slo__sro_n1620;
wire slo__n1187;
wire slo__n1188;
wire CLOCK_slo__sro_n1621;
wire CLOCK_slo__sro_n1622;
wire CLOCK_slo__sro_n1623;
wire CLOCK_slo__sro_n1624;
wire CLOCK_slo__sro_n1691;
wire CLOCK_slo__sro_n1692;
wire CLOCK_slo__sro_n1693;
wire CLOCK_slo__sro_n1694;
wire CLOCK_slo__sro_n1727;
wire CLOCK_slo__sro_n1728;
wire CLOCK_slo__sro_n1729;
wire CLOCK_slo__sro_n1730;
wire CLOCK_slo__sro_n1731;
wire CLOCK_slo__sro_n1746;
wire CLOCK_slo__sro_n1747;
wire CLOCK_slo__sro_n1748;
wire CLOCK_slo__sro_n1749;
wire CLOCK_slo__sro_n1759;
wire CLOCK_slo__sro_n1760;
wire slo__sro_n1535;
wire slo__sro_n1536;
wire slo__sro_n1537;
wire slo__sro_n1538;
wire slo__sro_n1539;
wire CLOCK_slo__mro_n1792;
wire CLOCK_slo__sro_n1786;


INV_X1 i_36 (.ZN (n_34), .A (p_0[30]));
INV_X2 i_35 (.ZN (n_33), .A (p_1[30]));
INV_X2 i_34 (.ZN (n_32), .A (n_30));
NAND2_X1 slo__sro_c635 (.ZN (slo__sro_n841), .A1 (p_1[18]), .A2 (p_0[18]));
XOR2_X2 i_32 (.Z (p_2[31]), .A (p_0[31]), .B (n_31));
OAI22_X1 i_31 (.ZN (n_0), .A1 (n_34), .A2 (p_1[30]), .B1 (n_33), .B2 (p_0[30]));
XNOR2_X1 i_0 (.ZN (p_2[30]), .A (n_32), .B (n_0));
INV_X1 CLOCK_slo__sro_c1311 (.ZN (CLOCK_slo__sro_n1694), .A (slo__sro_n271));
FA_X1 i_29 (.CO (n_29), .S (p_2[28]), .A (p_0[28]), .B (p_1[28]), .CI (n_28));
INV_X1 CLOCK_slo__sro_c1241 (.ZN (CLOCK_slo__sro_n1624), .A (slo__sro_n254));
FA_X1 i_27 (.CO (n_27), .S (p_2[26]), .A (p_0[26]), .B (p_1[26]), .CI (n_26));
FA_X1 i_26 (.CO (n_26), .S (p_2[25]), .A (p_0[25]), .B (p_1[25]), .CI (n_25));
FA_X1 i_25 (.CO (n_25), .S (p_2[24]), .A (p_0[24]), .B (p_1[24]), .CI (n_24));
FA_X1 i_24 (.CO (n_24), .S (p_2[23]), .A (p_0[23]), .B (p_1[23]), .CI (CLOCK_slo__sro_n1728));
INV_X1 CLOCK_slo__sro_c1362 (.ZN (CLOCK_slo__sro_n1749), .A (n_9));
FA_X1 i_22 (.CO (n_22), .S (p_2[21]), .A (p_0[21]), .B (p_1[21]), .CI (n_21));
INV_X1 CLOCK_slo__sro_c1346 (.ZN (CLOCK_slo__sro_n1731), .A (n_22));
INV_X1 slo__sro_c442 (.ZN (slo__sro_n594), .A (n_34));
XNOR2_X1 slo__sro_c783 (.ZN (slo__sro_n1026), .A (p_1[27]), .B (p_0[27]));
XNOR2_X1 slo__sro_c784 (.ZN (p_2[27]), .A (slo__sro_n1026), .B (n_27));
INV_X1 slo__sro_c68 (.ZN (slo__sro_n129), .A (p_1[2]));
INV_X1 CLOCK_slo__sro_c1255 (.ZN (CLOCK_slo__sro_n1637), .A (slo__sro_n590));
INV_X1 slo__sro_c202 (.ZN (slo__sro_n274), .A (slo__sro_n839));
INV_X1 slo__sro_c41 (.ZN (slo__sro_n104), .A (CLOCK_slo__sro_n1621));
INV_X2 slo__sro_c311 (.ZN (slo__sro_n391), .A (n_29));
FA_X1 i_12 (.CO (n_12), .S (p_2[11]), .A (p_0[11]), .B (p_1[11]), .CI (slo__sro_n344));
XNOR2_X1 slo__sro_c316 (.ZN (p_2[29]), .A (n_29), .B (slo__sro_n388));
CLKBUF_X1 spw__L1_c1_c2018 (.Z (spw_n2396), .A (p_1[30]));
FA_X1 i_9 (.CO (n_9), .S (p_2[8]), .A (p_0[8]), .B (p_1[8]), .CI (n_8));
FA_X1 i_8 (.CO (n_8), .S (p_2[7]), .A (p_0[7]), .B (p_1[7]), .CI (n_7));
FA_X1 i_7 (.CO (n_7), .S (p_2[6]), .A (p_0[6]), .B (p_1[6]), .CI (slo__sro_n1536));
XNOR2_X1 CLOCK_slo__mro_c1408 (.ZN (p_2[2]), .A (CLOCK_slo__mro_n1792), .B (n_2));
FA_X1 i_5 (.CO (n_5), .S (p_2[4]), .A (p_0[4]), .B (p_1[4]), .CI (CLOCK_slo__sro_n1760));
XNOR2_X1 CLOCK_slo__mro_c1407 (.ZN (CLOCK_slo__mro_n1792), .A (p_1[2]), .B (p_0[2]));
NAND2_X1 slo__sro_c203 (.ZN (slo__sro_n273), .A1 (p_1[19]), .A2 (p_0[19]));
FA_X1 i_2 (.CO (n_2), .S (p_2[1]), .A (p_0[1]), .B (p_1[1]), .CI (n_1));
HA_X1 i_1 (.CO (n_1), .S (p_2[0]), .A (p_0[0]), .B (p_1[0]));
NAND2_X1 CLOCK_slo__sro_c1257 (.ZN (CLOCK_slo__sro_n1635), .A1 (CLOCK_slo__sro_n1636), .A2 (CLOCK_slo__sro_n1637));
NAND2_X1 slo__sro_c189 (.ZN (slo__sro_n256), .A1 (p_1[14]), .A2 (p_0[14]));
NOR2_X1 slo__sro_c190 (.ZN (slo__sro_n255), .A1 (p_1[14]), .A2 (p_0[14]));
OAI21_X2 slo__sro_c191 (.ZN (slo__sro_n254), .A (slo__sro_n256), .B1 (slo__n1188), .B2 (slo__sro_n255));
XNOR2_X2 slo__sro_c192 (.ZN (slo__sro_n253), .A (p_1[14]), .B (p_0[14]));
XNOR2_X1 slo__sro_c193 (.ZN (p_2[14]), .A (slo__n1187), .B (slo__sro_n253));
INV_X1 slo__sro_c14 (.ZN (slo__sro_n76), .A (slo__sro_n302));
NAND2_X1 slo__sro_c15 (.ZN (slo__sro_n75), .A1 (p_1[13]), .A2 (p_0[13]));
NOR2_X1 slo__sro_c16 (.ZN (slo__sro_n74), .A1 (p_1[13]), .A2 (p_0[13]));
OAI21_X1 slo__sro_c17 (.ZN (n_14), .A (slo__sro_n75), .B1 (slo__sro_n74), .B2 (slo__sro_n76));
XNOR2_X1 slo__sro_c18 (.ZN (slo__sro_n73), .A (p_1[13]), .B (p_0[13]));
XNOR2_X1 slo__sro_c19 (.ZN (p_2[13]), .A (slo__sro_n73), .B (slo__sro_n302));
NAND2_X1 slo__sro_c42 (.ZN (slo__sro_n103), .A1 (p_1[16]), .A2 (p_0[16]));
NOR2_X1 slo__sro_c43 (.ZN (slo__sro_n102), .A1 (p_1[16]), .A2 (p_0[16]));
OAI21_X2 slo__sro_c44 (.ZN (n_17), .A (slo__sro_n103), .B1 (slo__sro_n104), .B2 (slo__sro_n102));
XNOR2_X1 slo__sro_c45 (.ZN (slo__sro_n101), .A (p_1[16]), .B (p_0[16]));
XNOR2_X1 slo__sro_c46 (.ZN (p_2[16]), .A (slo__sro_n101), .B (CLOCK_slo__sro_n1621));
NAND2_X1 slo__sro_c69 (.ZN (slo__sro_n128), .A1 (n_2), .A2 (p_0[2]));
NOR2_X2 slo__sro_c70 (.ZN (slo__sro_n127), .A1 (n_2), .A2 (p_0[2]));
OAI21_X1 slo__sro_c71 (.ZN (n_3), .A (slo__sro_n128), .B1 (slo__sro_n129), .B2 (slo__sro_n127));
NOR2_X1 slo__sro_c204 (.ZN (slo__sro_n272), .A1 (p_1[19]), .A2 (p_0[19]));
OAI21_X2 slo__sro_c205 (.ZN (slo__sro_n271), .A (slo__sro_n273), .B1 (slo__sro_n274), .B2 (slo__sro_n272));
XNOR2_X2 slo__sro_c206 (.ZN (slo__sro_n270), .A (p_1[19]), .B (p_0[19]));
XNOR2_X2 slo__sro_c207 (.ZN (p_2[19]), .A (slo__sro_n270), .B (slo__sro_n839));
INV_X1 slo__sro_c443 (.ZN (slo__sro_n593), .A (spw_n2396));
INV_X1 slo__sro_c444 (.ZN (slo__sro_n592), .A (n_33));
INV_X1 slo__sro_c445 (.ZN (slo__sro_n591), .A (p_0[30]));
NAND2_X1 slo__sro_c446 (.ZN (slo__sro_n590), .A1 (slo__sro_n592), .A2 (slo__sro_n591));
NAND2_X1 slo__sro_c447 (.ZN (slo__sro_n589), .A1 (slo__sro_n593), .A2 (slo__sro_n594));
INV_X1 slo__sro_c231 (.ZN (slo__sro_n305), .A (n_12));
NAND2_X1 slo__sro_c232 (.ZN (slo__sro_n304), .A1 (p_1[12]), .A2 (p_0[12]));
NOR2_X1 slo__sro_c233 (.ZN (slo__sro_n303), .A1 (p_1[12]), .A2 (p_0[12]));
OAI21_X2 slo__sro_c234 (.ZN (slo__sro_n302), .A (slo__sro_n304), .B1 (slo__sro_n305), .B2 (slo__sro_n303));
XNOR2_X1 slo__sro_c235 (.ZN (slo__sro_n301), .A (p_1[12]), .B (p_0[12]));
XNOR2_X2 slo__sro_c236 (.ZN (p_2[12]), .A (n_12), .B (slo__sro_n301));
NAND2_X1 slo__sro_c312 (.ZN (slo__sro_n390), .A1 (p_1[29]), .A2 (p_0[29]));
NOR2_X1 slo__sro_c313 (.ZN (slo__sro_n389), .A1 (p_1[29]), .A2 (p_0[29]));
OAI21_X2 slo__sro_c314 (.ZN (n_30), .A (slo__sro_n390), .B1 (slo__sro_n391), .B2 (slo__sro_n389));
XNOR2_X1 slo__sro_c315 (.ZN (slo__sro_n388), .A (p_1[29]), .B (p_0[29]));
INV_X1 slo__sro_c271 (.ZN (slo__sro_n347), .A (n_10));
NAND2_X1 slo__sro_c272 (.ZN (slo__sro_n346), .A1 (p_1[10]), .A2 (p_0[10]));
NOR2_X1 slo__sro_c273 (.ZN (slo__sro_n345), .A1 (p_1[10]), .A2 (p_0[10]));
OAI21_X1 slo__sro_c274 (.ZN (slo__sro_n344), .A (slo__sro_n346), .B1 (slo__sro_n347), .B2 (slo__sro_n345));
XNOR2_X1 slo__sro_c275 (.ZN (slo__sro_n343), .A (p_1[10]), .B (p_0[10]));
XNOR2_X1 slo__sro_c276 (.ZN (p_2[10]), .A (slo__sro_n343), .B (n_10));
OAI21_X1 slo__sro_c636 (.ZN (slo__sro_n840), .A (slo__sro_n721), .B1 (p_1[18]), .B2 (p_0[18]));
NAND2_X2 slo__sro_c637 (.ZN (slo__sro_n839), .A1 (slo__sro_n840), .A2 (slo__sro_n841));
XNOR2_X2 slo__sro_c638 (.ZN (slo__sro_n838), .A (p_1[18]), .B (p_0[18]));
XNOR2_X2 slo__sro_c639 (.ZN (p_2[18]), .A (slo__sro_n838), .B (slo__sro_n721));
NAND2_X1 slo__sro_c567 (.ZN (slo__sro_n723), .A1 (p_1[17]), .A2 (p_0[17]));
INV_X2 slo__sro_c779 (.ZN (slo__sro_n1029), .A (n_27));
NAND2_X2 slo__sro_c569 (.ZN (slo__sro_n721), .A1 (slo__sro_n1014), .A2 (slo__sro_n723));
XNOR2_X1 slo__sro_c570 (.ZN (slo__sro_n720), .A (p_1[17]), .B (p_0[17]));
XNOR2_X2 slo__sro_c571 (.ZN (p_2[17]), .A (slo__sro_n720), .B (n_17));
INV_X1 slo__sro_c769 (.ZN (slo__sro_n1017), .A (p_1[17]));
INV_X1 slo__sro_c770 (.ZN (slo__sro_n1016), .A (p_0[17]));
NAND2_X1 slo__sro_c771 (.ZN (slo__sro_n1015), .A1 (slo__sro_n1017), .A2 (slo__sro_n1016));
NAND2_X1 slo__sro_c772 (.ZN (slo__sro_n1014), .A1 (n_17), .A2 (slo__sro_n1015));
NAND2_X1 slo__sro_c780 (.ZN (slo__sro_n1028), .A1 (p_0[27]), .A2 (p_1[27]));
NOR2_X2 slo__sro_c781 (.ZN (slo__sro_n1027), .A1 (p_1[27]), .A2 (p_0[27]));
OAI21_X2 slo__sro_c782 (.ZN (n_28), .A (slo__sro_n1028), .B1 (slo__sro_n1029), .B2 (slo__sro_n1027));
NAND2_X1 CLOCK_slo__sro_c1242 (.ZN (CLOCK_slo__sro_n1623), .A1 (p_1[15]), .A2 (p_0[15]));
OAI21_X1 CLOCK_slo__sro_c1258 (.ZN (n_31), .A (CLOCK_slo__sro_n1635), .B1 (n_32), .B2 (slo__sro_n589));
CLKBUF_X1 slo__L1_c909 (.Z (slo__n1187), .A (n_14));
INV_X1 slo__L1_c910 (.ZN (slo__n1188), .A (n_14));
NOR2_X1 CLOCK_slo__sro_c1243 (.ZN (CLOCK_slo__sro_n1622), .A1 (p_1[15]), .A2 (p_0[15]));
OAI21_X2 CLOCK_slo__sro_c1244 (.ZN (CLOCK_slo__sro_n1621), .A (CLOCK_slo__sro_n1623)
    , .B1 (CLOCK_slo__sro_n1624), .B2 (CLOCK_slo__sro_n1622));
XNOR2_X1 CLOCK_slo__sro_c1245 (.ZN (CLOCK_slo__sro_n1620), .A (p_1[15]), .B (p_0[15]));
XNOR2_X1 CLOCK_slo__sro_c1246 (.ZN (p_2[15]), .A (CLOCK_slo__sro_n1620), .B (slo__sro_n254));
INV_X1 CLOCK_slo__sro_c1256 (.ZN (CLOCK_slo__sro_n1636), .A (n_30));
NAND2_X1 CLOCK_slo__sro_c1312 (.ZN (CLOCK_slo__sro_n1693), .A1 (p_1[20]), .A2 (p_0[20]));
NOR2_X1 CLOCK_slo__sro_c1313 (.ZN (CLOCK_slo__sro_n1692), .A1 (p_1[20]), .A2 (p_0[20]));
OAI21_X1 CLOCK_slo__sro_c1314 (.ZN (n_21), .A (CLOCK_slo__sro_n1693), .B1 (CLOCK_slo__sro_n1694), .B2 (CLOCK_slo__sro_n1692));
XNOR2_X1 CLOCK_slo__sro_c1315 (.ZN (CLOCK_slo__sro_n1691), .A (p_1[20]), .B (p_0[20]));
XNOR2_X1 CLOCK_slo__sro_c1316 (.ZN (p_2[20]), .A (CLOCK_slo__sro_n1691), .B (slo__sro_n271));
NAND2_X1 CLOCK_slo__sro_c1347 (.ZN (CLOCK_slo__sro_n1730), .A1 (p_1[22]), .A2 (p_0[22]));
NOR2_X2 CLOCK_slo__sro_c1348 (.ZN (CLOCK_slo__sro_n1729), .A1 (p_1[22]), .A2 (p_0[22]));
OAI21_X1 CLOCK_slo__sro_c1349 (.ZN (CLOCK_slo__sro_n1728), .A (CLOCK_slo__sro_n1730)
    , .B1 (CLOCK_slo__sro_n1731), .B2 (CLOCK_slo__sro_n1729));
XNOR2_X1 CLOCK_slo__sro_c1350 (.ZN (CLOCK_slo__sro_n1727), .A (p_1[22]), .B (p_0[22]));
XNOR2_X1 CLOCK_slo__sro_c1351 (.ZN (p_2[22]), .A (CLOCK_slo__sro_n1727), .B (n_22));
NAND2_X1 CLOCK_slo__sro_c1363 (.ZN (CLOCK_slo__sro_n1748), .A1 (p_1[9]), .A2 (p_0[9]));
NOR2_X1 CLOCK_slo__sro_c1364 (.ZN (CLOCK_slo__sro_n1747), .A1 (p_1[9]), .A2 (p_0[9]));
OAI21_X2 CLOCK_slo__sro_c1365 (.ZN (n_10), .A (CLOCK_slo__sro_n1748), .B1 (CLOCK_slo__sro_n1749), .B2 (CLOCK_slo__sro_n1747));
XNOR2_X1 CLOCK_slo__sro_c1366 (.ZN (CLOCK_slo__sro_n1746), .A (p_1[9]), .B (p_0[9]));
XNOR2_X1 CLOCK_slo__sro_c1367 (.ZN (p_2[9]), .A (n_9), .B (CLOCK_slo__sro_n1746));
NAND2_X1 CLOCK_slo__sro_c1377 (.ZN (CLOCK_slo__sro_n1762), .A1 (p_1[3]), .A2 (p_0[3]));
NAND2_X1 CLOCK_slo__sro_c1379 (.ZN (CLOCK_slo__sro_n1760), .A1 (CLOCK_slo__sro_n1786), .A2 (CLOCK_slo__sro_n1762));
XNOR2_X1 CLOCK_slo__sro_c1380 (.ZN (CLOCK_slo__sro_n1759), .A (n_3), .B (p_0[3]));
XNOR2_X1 CLOCK_slo__sro_c1381 (.ZN (p_2[3]), .A (CLOCK_slo__sro_n1759), .B (p_1[3]));
INV_X1 slo__sro_c1188 (.ZN (slo__sro_n1539), .A (n_5));
NAND2_X1 slo__sro_c1189 (.ZN (slo__sro_n1538), .A1 (p_1[5]), .A2 (p_0[5]));
NOR2_X1 slo__sro_c1190 (.ZN (slo__sro_n1537), .A1 (p_1[5]), .A2 (p_0[5]));
OAI21_X1 slo__sro_c1191 (.ZN (slo__sro_n1536), .A (slo__sro_n1538), .B1 (slo__sro_n1539), .B2 (slo__sro_n1537));
XNOR2_X2 slo__sro_c1192 (.ZN (slo__sro_n1535), .A (p_1[5]), .B (p_0[5]));
XNOR2_X1 slo__sro_c1193 (.ZN (p_2[5]), .A (slo__sro_n1535), .B (n_5));
OAI21_X1 CLOCK_slo__sro_c1403 (.ZN (CLOCK_slo__sro_n1786), .A (n_3), .B1 (p_1[3]), .B2 (p_0[3]));

endmodule //datapath__0_232

module datapath__0_231 (Multiplier, p_0, p_1);

output [31:0] p_1;
input [31:0] Multiplier;
input [31:0] p_0;
wire n_1;
wire n_2;
wire n_3;
wire n_4;
wire n_5;
wire n_6;
wire n_7;
wire n_8;
wire n_10;
wire n_11;
wire n_12;
wire n_13;
wire n_16;
wire n_18;
wire n_19;
wire n_21;
wire n_22;
wire n_23;
wire n_25;
wire n_27;
wire n_29;
wire n_30;
wire n_32;
wire n_34;
wire n_33;
wire slo__sro_n59;
wire slo__sro_n60;
wire slo__sro_n61;
wire slo__sro_n62;
wire slo__sro_n72;
wire slo__sro_n73;
wire slo__sro_n74;
wire slo__sro_n75;
wire slo__sro_n76;
wire slo__sro_n89;
wire slo__sro_n90;
wire slo__sro_n91;
wire slo__sro_n92;
wire slo__sro_n102;
wire slo__sro_n103;
wire slo__sro_n104;
wire slo__sro_n105;
wire slo__sro_n106;
wire slo__sro_n119;
wire slo__sro_n120;
wire slo__sro_n121;
wire slo__sro_n122;
wire slo__sro_n123;
wire slo__sro_n138;
wire slo__sro_n139;
wire slo__sro_n140;
wire slo__sro_n151;
wire slo__sro_n152;
wire slo__sro_n153;
wire slo__sro_n154;
wire slo__sro_n166;
wire slo__sro_n167;
wire slo__sro_n168;
wire slo__sro_n169;
wire slo__sro_n844;
wire CLOCK_slo__sro_n1021;
wire slo__sro_n180;
wire slo__sro_n181;
wire slo__sro_n182;
wire slo__sro_n183;
wire slo__sro_n198;
wire slo__sro_n199;
wire slo__sro_n200;
wire slo__sro_n201;
wire slo__sro_n202;
wire slo__sro_n217;
wire slo__sro_n218;
wire slo__sro_n219;
wire slo__sro_n220;
wire slo__sro_n221;
wire slo__sro_n234;
wire slo__sro_n235;
wire slo__sro_n236;
wire slo__sro_n237;
wire slo__sro_n238;
wire slo__sro_n251;
wire slo__sro_n252;
wire slo__sro_n253;
wire slo__sro_n260;
wire slo__sro_n261;
wire slo__sro_n262;
wire slo__sro_n263;
wire slo__sro_n264;
wire slo__sro_n727;
wire slo__sro_n728;
wire slo__sro_n729;
wire slo__sro_n730;
wire CLOCK_slo__sro_n1022;
wire CLOCK_slo__sro_n1023;
wire CLOCK_slo__sro_n1047;
wire slo__sro_n871;
wire CLOCK_slo__sro_n1048;
wire CLOCK_slo__sro_n1049;
wire CLOCK_slo__sro_n1050;
wire CLOCK_slo__sro_n1108;
wire CLOCK_slo__sro_n1109;
wire CLOCK_slo__sro_n1110;
wire CLOCK_slo__sro_n1111;
wire CLOCK_slo__sro_n1112;
wire CLOCK_slo__sro_n1142;
wire CLOCK_slo__sro_n1143;
wire CLOCK_slo__sro_n1144;
wire CLOCK_slo__sro_n1145;
wire CLOCK_slo__sro_n1157;
wire CLOCK_slo__sro_n1158;
wire CLOCK_slo__sro_n1159;
wire CLOCK_slo__sro_n1160;
wire CLOCK_slo__sro_n1371;
wire CLOCK_slo__sro_n1372;
wire CLOCK_slo__sro_n1373;


INV_X1 i_36 (.ZN (n_34), .A (Multiplier[30]));
INV_X2 i_35 (.ZN (n_33), .A (p_0[30]));
INV_X2 i_34 (.ZN (n_32), .A (n_30));
XOR2_X1 i_32 (.Z (p_1[31]), .A (slo__sro_n260), .B (Multiplier[31]));
XNOR2_X2 i_0 (.ZN (p_1[30]), .A (n_32), .B (slo__sro_n871));
INV_X1 CLOCK_slo__sro_c728 (.ZN (CLOCK_slo__sro_n1112), .A (n_23));
FA_X1 i_29 (.CO (n_29), .S (p_1[28]), .A (Multiplier[28]), .B (p_0[28]), .CI (slo__sro_n235));
NAND2_X1 slo__sro_c175 (.ZN (slo__sro_n253), .A1 (n_10), .A2 (Multiplier[10]));
FA_X1 i_27 (.CO (n_27), .S (p_1[26]), .A (Multiplier[26]), .B (p_0[26]), .CI (slo__sro_n103));
INV_X1 slo__sro_c59 (.ZN (slo__sro_n123), .A (n_19));
INV_X1 slo__sro_c87 (.ZN (slo__sro_n154), .A (n_22));
INV_X1 CLOCK_slo__sro_c765 (.ZN (CLOCK_slo__sro_n1145), .A (n_11));
INV_X4 slo__sro_c101 (.ZN (slo__sro_n169), .A (slo__sro_n199));
FA_X1 i_22 (.CO (n_22), .S (p_1[21]), .A (Multiplier[21]), .B (p_0[21]), .CI (n_21));
FA_X1 i_21 (.CO (n_21), .S (p_1[20]), .A (Multiplier[20]), .B (p_0[20]), .CI (slo__sro_n120));
NAND2_X1 slo__sro_c75 (.ZN (slo__sro_n140), .A1 (p_0[24]), .A2 (Multiplier[24]));
FA_X1 i_19 (.CO (n_19), .S (p_1[18]), .A (Multiplier[18]), .B (p_0[18]), .CI (n_18));
XNOR2_X2 slo__sro_c533 (.ZN (p_1[13]), .A (slo__sro_n844), .B (n_13));
INV_X1 slo__sro_c31 (.ZN (slo__sro_n92), .A (n_2));
INV_X2 slo__sro_c17 (.ZN (slo__sro_n76), .A (p_0[16]));
INV_X1 slo__sro_c161 (.ZN (slo__sro_n238), .A (n_27));
INV_X1 slo__sro_c131 (.ZN (slo__sro_n202), .A (n_8));
FA_X1 i_13 (.CO (n_13), .S (p_1[12]), .A (Multiplier[12]), .B (p_0[12]), .CI (n_12));
NAND2_X1 CLOCK_slo__sro_c781 (.ZN (CLOCK_slo__sro_n1160), .A1 (p_0[4]), .A2 (Multiplier[4]));
INV_X1 slo__sro_c187 (.ZN (slo__sro_n264), .A (n_30));
INV_X1 slo__sro_c115 (.ZN (slo__sro_n183), .A (n_13));
INV_X1 slo__sro_c147 (.ZN (slo__sro_n221), .A (p_0[14]));
FA_X1 i_8 (.CO (n_8), .S (p_1[7]), .A (Multiplier[7]), .B (p_0[7]), .CI (n_7));
FA_X1 i_7 (.CO (n_7), .S (p_1[6]), .A (Multiplier[6]), .B (p_0[6]), .CI (n_6));
FA_X1 i_6 (.CO (n_6), .S (p_1[5]), .A (Multiplier[5]), .B (p_0[5]), .CI (n_5));
INV_X1 CLOCK_slo__sro_c668 (.ZN (CLOCK_slo__sro_n1050), .A (n_29));
INV_X1 slo__sro_c45 (.ZN (slo__sro_n106), .A (n_25));
HA_X1 i_1 (.CO (n_1), .S (p_1[0]), .A (Multiplier[0]), .B (p_0[0]));
INV_X1 slo__sro_c3 (.ZN (slo__sro_n62), .A (slo__sro_n218));
NAND2_X1 slo__sro_c4 (.ZN (slo__sro_n61), .A1 (p_0[15]), .A2 (Multiplier[15]));
NOR2_X2 slo__sro_c5 (.ZN (slo__sro_n60), .A1 (p_0[15]), .A2 (Multiplier[15]));
OAI21_X2 slo__sro_c6 (.ZN (n_16), .A (slo__sro_n61), .B1 (slo__sro_n62), .B2 (slo__sro_n60));
XNOR2_X1 slo__sro_c7 (.ZN (slo__sro_n59), .A (p_0[15]), .B (Multiplier[15]));
XNOR2_X1 slo__sro_c8 (.ZN (p_1[15]), .A (slo__sro_n59), .B (slo__sro_n218));
NAND2_X1 slo__sro_c18 (.ZN (slo__sro_n75), .A1 (n_16), .A2 (Multiplier[16]));
NOR2_X2 slo__sro_c19 (.ZN (slo__sro_n74), .A1 (n_16), .A2 (Multiplier[16]));
OAI21_X2 slo__sro_c20 (.ZN (slo__sro_n73), .A (slo__sro_n75), .B1 (slo__sro_n74), .B2 (slo__sro_n76));
XNOR2_X1 slo__sro_c21 (.ZN (slo__sro_n72), .A (n_16), .B (Multiplier[16]));
XNOR2_X2 slo__sro_c22 (.ZN (p_1[16]), .A (slo__sro_n72), .B (p_0[16]));
NAND2_X1 slo__sro_c32 (.ZN (slo__sro_n91), .A1 (p_0[2]), .A2 (Multiplier[2]));
NOR2_X2 slo__sro_c33 (.ZN (slo__sro_n90), .A1 (p_0[2]), .A2 (Multiplier[2]));
OAI21_X2 slo__sro_c34 (.ZN (n_3), .A (slo__sro_n91), .B1 (slo__sro_n92), .B2 (slo__sro_n90));
XNOR2_X2 slo__sro_c35 (.ZN (slo__sro_n89), .A (p_0[2]), .B (Multiplier[2]));
XNOR2_X2 slo__sro_c36 (.ZN (p_1[2]), .A (slo__sro_n89), .B (n_2));
NAND2_X1 slo__sro_c46 (.ZN (slo__sro_n105), .A1 (p_0[25]), .A2 (Multiplier[25]));
NOR2_X2 slo__sro_c47 (.ZN (slo__sro_n104), .A1 (p_0[25]), .A2 (Multiplier[25]));
OAI21_X1 slo__sro_c48 (.ZN (slo__sro_n103), .A (slo__sro_n105), .B1 (slo__sro_n104), .B2 (slo__sro_n106));
XNOR2_X2 slo__sro_c49 (.ZN (slo__sro_n102), .A (p_0[25]), .B (Multiplier[25]));
XNOR2_X2 slo__sro_c50 (.ZN (p_1[25]), .A (slo__sro_n102), .B (n_25));
NAND2_X1 slo__sro_c60 (.ZN (slo__sro_n122), .A1 (p_0[19]), .A2 (Multiplier[19]));
NOR2_X1 slo__sro_c61 (.ZN (slo__sro_n121), .A1 (p_0[19]), .A2 (Multiplier[19]));
NAND2_X1 CLOCK_slo__sro_c640 (.ZN (CLOCK_slo__sro_n1023), .A1 (p_0[3]), .A2 (Multiplier[3]));
XNOR2_X1 slo__sro_c63 (.ZN (slo__sro_n119), .A (p_0[19]), .B (Multiplier[19]));
XNOR2_X2 slo__sro_c64 (.ZN (p_1[19]), .A (n_19), .B (slo__sro_n119));
OAI21_X1 slo__sro_c76 (.ZN (slo__sro_n139), .A (CLOCK_slo__sro_n1109), .B1 (p_0[24]), .B2 (Multiplier[24]));
NAND2_X1 slo__sro_c77 (.ZN (n_25), .A1 (slo__sro_n140), .A2 (slo__sro_n139));
XNOR2_X2 slo__sro_c78 (.ZN (slo__sro_n138), .A (p_0[24]), .B (Multiplier[24]));
XNOR2_X1 slo__sro_c79 (.ZN (p_1[24]), .A (slo__sro_n138), .B (CLOCK_slo__sro_n1109));
NAND2_X1 slo__sro_c88 (.ZN (slo__sro_n153), .A1 (p_0[22]), .A2 (Multiplier[22]));
NOR2_X1 slo__sro_c89 (.ZN (slo__sro_n152), .A1 (p_0[22]), .A2 (Multiplier[22]));
OAI21_X2 slo__sro_c90 (.ZN (n_23), .A (slo__sro_n153), .B1 (slo__sro_n154), .B2 (slo__sro_n152));
XNOR2_X1 slo__sro_c91 (.ZN (slo__sro_n151), .A (p_0[22]), .B (Multiplier[22]));
XNOR2_X1 slo__sro_c92 (.ZN (p_1[22]), .A (n_22), .B (slo__sro_n151));
NAND2_X1 slo__sro_c102 (.ZN (slo__sro_n168), .A1 (p_0[9]), .A2 (Multiplier[9]));
NOR2_X1 slo__sro_c103 (.ZN (slo__sro_n167), .A1 (p_0[9]), .A2 (Multiplier[9]));
OAI21_X2 slo__sro_c104 (.ZN (n_10), .A (slo__sro_n168), .B1 (slo__sro_n167), .B2 (slo__sro_n169));
XNOR2_X1 slo__sro_c105 (.ZN (slo__sro_n166), .A (p_0[9]), .B (Multiplier[9]));
XNOR2_X1 slo__sro_c106 (.ZN (p_1[9]), .A (slo__sro_n166), .B (slo__sro_n199));
NAND2_X1 slo__sro_c116 (.ZN (slo__sro_n182), .A1 (p_0[13]), .A2 (Multiplier[13]));
NOR2_X1 slo__sro_c117 (.ZN (slo__sro_n181), .A1 (p_0[13]), .A2 (Multiplier[13]));
OAI21_X2 slo__sro_c118 (.ZN (slo__sro_n180), .A (slo__sro_n182), .B1 (slo__sro_n183), .B2 (slo__sro_n181));
OAI21_X2 CLOCK_slo__sro_c641 (.ZN (CLOCK_slo__sro_n1022), .A (n_3), .B1 (p_0[3]), .B2 (Multiplier[3]));
XNOR2_X2 slo__sro_c542 (.ZN (slo__sro_n844), .A (p_0[13]), .B (Multiplier[13]));
NAND2_X1 slo__sro_c132 (.ZN (slo__sro_n201), .A1 (p_0[8]), .A2 (Multiplier[8]));
NOR2_X1 slo__sro_c133 (.ZN (slo__sro_n200), .A1 (p_0[8]), .A2 (Multiplier[8]));
OAI21_X4 slo__sro_c134 (.ZN (slo__sro_n199), .A (slo__sro_n201), .B1 (slo__sro_n200), .B2 (slo__sro_n202));
XNOR2_X1 slo__sro_c135 (.ZN (slo__sro_n198), .A (p_0[8]), .B (Multiplier[8]));
XNOR2_X1 slo__sro_c136 (.ZN (p_1[8]), .A (slo__sro_n198), .B (n_8));
NAND2_X1 slo__sro_c148 (.ZN (slo__sro_n220), .A1 (slo__sro_n180), .A2 (Multiplier[14]));
NOR2_X2 slo__sro_c149 (.ZN (slo__sro_n219), .A1 (slo__sro_n180), .A2 (Multiplier[14]));
NAND2_X1 CLOCK_slo__sro_c975 (.ZN (n_2), .A1 (CLOCK_slo__sro_n1372), .A2 (CLOCK_slo__sro_n1373));
XNOR2_X1 slo__sro_c151 (.ZN (slo__sro_n217), .A (slo__sro_n180), .B (Multiplier[14]));
XNOR2_X1 slo__sro_c152 (.ZN (p_1[14]), .A (slo__sro_n217), .B (p_0[14]));
NAND2_X1 slo__sro_c162 (.ZN (slo__sro_n237), .A1 (p_0[27]), .A2 (Multiplier[27]));
NOR2_X1 slo__sro_c163 (.ZN (slo__sro_n236), .A1 (p_0[27]), .A2 (Multiplier[27]));
OAI21_X1 slo__sro_c164 (.ZN (slo__sro_n235), .A (slo__sro_n237), .B1 (slo__sro_n236), .B2 (slo__sro_n238));
XNOR2_X1 slo__sro_c165 (.ZN (slo__sro_n234), .A (p_0[27]), .B (Multiplier[27]));
XNOR2_X1 slo__sro_c166 (.ZN (p_1[27]), .A (slo__sro_n234), .B (n_27));
OAI21_X1 slo__sro_c176 (.ZN (slo__sro_n252), .A (p_0[10]), .B1 (n_10), .B2 (Multiplier[10]));
NAND2_X1 slo__sro_c177 (.ZN (n_11), .A1 (slo__sro_n252), .A2 (slo__sro_n253));
XNOR2_X1 slo__sro_c178 (.ZN (slo__sro_n251), .A (n_10), .B (Multiplier[10]));
XNOR2_X1 slo__sro_c179 (.ZN (p_1[10]), .A (slo__sro_n251), .B (p_0[10]));
NOR2_X1 slo__sro_c188 (.ZN (slo__sro_n263), .A1 (n_33), .A2 (Multiplier[30]));
NAND2_X1 slo__sro_c189 (.ZN (slo__sro_n262), .A1 (slo__sro_n263), .A2 (slo__sro_n264));
OR2_X1 slo__sro_c190 (.ZN (slo__sro_n261), .A1 (p_0[30]), .A2 (n_34));
OAI21_X2 slo__sro_c191 (.ZN (slo__sro_n260), .A (slo__sro_n262), .B1 (n_32), .B2 (slo__sro_n261));
OAI21_X1 slo__sro_c562 (.ZN (slo__sro_n120), .A (slo__sro_n122), .B1 (slo__sro_n123), .B2 (slo__sro_n121));
NAND2_X1 slo__sro_c474 (.ZN (slo__sro_n730), .A1 (p_0[17]), .A2 (Multiplier[17]));
NAND2_X1 slo__sro_c475 (.ZN (slo__sro_n729), .A1 (slo__sro_n73), .A2 (Multiplier[17]));
NAND2_X2 slo__sro_c476 (.ZN (slo__sro_n728), .A1 (slo__sro_n73), .A2 (p_0[17]));
NAND3_X2 slo__sro_c477 (.ZN (n_18), .A1 (slo__sro_n729), .A2 (slo__sro_n728), .A3 (slo__sro_n730));
XNOR2_X1 slo__sro_c478 (.ZN (slo__sro_n727), .A (p_0[17]), .B (Multiplier[17]));
XNOR2_X1 slo__sro_c479 (.ZN (p_1[17]), .A (slo__sro_n727), .B (slo__sro_n73));
NAND2_X2 CLOCK_slo__sro_c642 (.ZN (n_4), .A1 (CLOCK_slo__sro_n1023), .A2 (CLOCK_slo__sro_n1022));
XNOR2_X1 CLOCK_slo__sro_c643 (.ZN (CLOCK_slo__sro_n1021), .A (n_3), .B (Multiplier[3]));
OAI22_X2 slo__sro_c558 (.ZN (slo__sro_n871), .A1 (n_33), .A2 (Multiplier[30]), .B1 (p_0[30]), .B2 (n_34));
XNOR2_X1 CLOCK_slo__sro_c644 (.ZN (p_1[3]), .A (CLOCK_slo__sro_n1021), .B (p_0[3]));
NAND2_X1 CLOCK_slo__sro_c669 (.ZN (CLOCK_slo__sro_n1049), .A1 (p_0[29]), .A2 (Multiplier[29]));
NOR2_X2 CLOCK_slo__sro_c670 (.ZN (CLOCK_slo__sro_n1048), .A1 (p_0[29]), .A2 (Multiplier[29]));
OAI21_X2 CLOCK_slo__sro_c671 (.ZN (n_30), .A (CLOCK_slo__sro_n1049), .B1 (CLOCK_slo__sro_n1050), .B2 (CLOCK_slo__sro_n1048));
XNOR2_X1 CLOCK_slo__sro_c672 (.ZN (CLOCK_slo__sro_n1047), .A (p_0[29]), .B (Multiplier[29]));
XNOR2_X1 CLOCK_slo__sro_c673 (.ZN (p_1[29]), .A (CLOCK_slo__sro_n1047), .B (n_29));
NAND2_X1 CLOCK_slo__sro_c729 (.ZN (CLOCK_slo__sro_n1111), .A1 (p_0[23]), .A2 (Multiplier[23]));
NOR2_X1 CLOCK_slo__sro_c730 (.ZN (CLOCK_slo__sro_n1110), .A1 (p_0[23]), .A2 (Multiplier[23]));
OAI21_X1 CLOCK_slo__sro_c731 (.ZN (CLOCK_slo__sro_n1109), .A (CLOCK_slo__sro_n1111)
    , .B1 (CLOCK_slo__sro_n1112), .B2 (CLOCK_slo__sro_n1110));
XNOR2_X1 CLOCK_slo__sro_c732 (.ZN (CLOCK_slo__sro_n1108), .A (p_0[23]), .B (Multiplier[23]));
XNOR2_X1 CLOCK_slo__sro_c733 (.ZN (p_1[23]), .A (CLOCK_slo__sro_n1108), .B (n_23));
NAND2_X1 CLOCK_slo__sro_c766 (.ZN (CLOCK_slo__sro_n1144), .A1 (p_0[11]), .A2 (Multiplier[11]));
NOR2_X1 CLOCK_slo__sro_c767 (.ZN (CLOCK_slo__sro_n1143), .A1 (p_0[11]), .A2 (Multiplier[11]));
OAI21_X1 CLOCK_slo__sro_c768 (.ZN (n_12), .A (CLOCK_slo__sro_n1144), .B1 (CLOCK_slo__sro_n1145), .B2 (CLOCK_slo__sro_n1143));
XNOR2_X1 CLOCK_slo__sro_c769 (.ZN (CLOCK_slo__sro_n1142), .A (p_0[11]), .B (Multiplier[11]));
XNOR2_X1 CLOCK_slo__sro_c770 (.ZN (p_1[11]), .A (CLOCK_slo__sro_n1142), .B (n_11));
NAND2_X1 CLOCK_slo__sro_c782 (.ZN (CLOCK_slo__sro_n1159), .A1 (n_4), .A2 (Multiplier[4]));
NAND2_X1 CLOCK_slo__sro_c783 (.ZN (CLOCK_slo__sro_n1158), .A1 (p_0[4]), .A2 (n_4));
NAND3_X1 CLOCK_slo__sro_c784 (.ZN (n_5), .A1 (CLOCK_slo__sro_n1160), .A2 (CLOCK_slo__sro_n1158), .A3 (CLOCK_slo__sro_n1159));
XNOR2_X2 CLOCK_slo__sro_c785 (.ZN (CLOCK_slo__sro_n1157), .A (n_4), .B (Multiplier[4]));
XNOR2_X2 CLOCK_slo__sro_c786 (.ZN (p_1[4]), .A (CLOCK_slo__sro_n1157), .B (p_0[4]));
NAND2_X1 CLOCK_slo__sro_c973 (.ZN (CLOCK_slo__sro_n1373), .A1 (n_1), .A2 (Multiplier[1]));
AOI22_X1 CLOCK_slo__sro_c974 (.ZN (CLOCK_slo__sro_n1372), .A1 (n_1), .A2 (p_0[1])
    , .B1 (p_0[1]), .B2 (Multiplier[1]));
OAI21_X2 CLOCK_slo__sro_c888 (.ZN (slo__sro_n218), .A (slo__sro_n220), .B1 (slo__sro_n219), .B2 (slo__sro_n221));
XNOR2_X1 CLOCK_slo__sro_c976 (.ZN (CLOCK_slo__sro_n1371), .A (p_0[1]), .B (Multiplier[1]));
XNOR2_X1 CLOCK_slo__sro_c977 (.ZN (p_1[1]), .A (CLOCK_slo__sro_n1371), .B (n_1));

endmodule //datapath__0_231

module datapath__0_227 (p_1_22_PP_5, p_0, p_1, p_2);

output [31:0] p_2;
input [31:0] p_0;
input [31:0] p_1;
input p_1_22_PP_5;
wire CLOCK_slo__sro_n1768;
wire CLOCK_slo__sro_n1381;
wire n_1;
wire n_2;
wire n_4;
wire n_5;
wire n_6;
wire n_7;
wire slo__sro_n237;
wire n_9;
wire n_10;
wire n_12;
wire n_13;
wire n_14;
wire n_15;
wire n_16;
wire slo__sro_n610;
wire n_19;
wire n_20;
wire n_21;
wire n_25;
wire n_26;
wire n_29;
wire n_30;
wire n_32;
wire n_0;
wire n_34;
wire n_33;
wire slo__sro_n63;
wire slo__sro_n64;
wire slo__sro_n65;
wire slo__sro_n66;
wire slo__sro_n76;
wire slo__sro_n77;
wire slo__sro_n78;
wire slo__sro_n79;
wire slo__sro_n80;
wire slo__sro_n93;
wire slo__sro_n94;
wire slo__sro_n95;
wire slo__sro_n96;
wire slo__sro_n97;
wire slo__sro_n112;
wire slo__sro_n113;
wire slo__sro_n114;
wire slo__sro_n115;
wire CLOCK_slo__sro_n1431;
wire slo__sro_n143;
wire slo__sro_n144;
wire CLOCK_slo__sro_n1382;
wire slo__sro_n146;
wire slo__sro_n220;
wire CLOCK_slo__mro_n1314;
wire slo__sro_n222;
wire slo__sro_n223;
wire slo__sro_n171;
wire slo__sro_n172;
wire slo__sro_n173;
wire slo__sro_n174;
wire slo__sro_n224;
wire slo__sro_n225;
wire slo__sro_n238;
wire slo__sro_n239;
wire slo__sro_n240;
wire slo__sro_n241;
wire CLOCK_slo__sro_n1331;
wire slo__n265;
wire slo__sro_n609;
wire slo__sro_n309;
wire slo__sro_n310;
wire slo__sro_n311;
wire slo__sro_n312;
wire slo__sro_n362;
wire slo__sro_n363;
wire slo__sro_n364;
wire slo__sro_n365;
wire slo__sro_n366;
wire slo__sro_n439;
wire slo__sro_n440;
wire slo__sro_n441;
wire slo__sro_n442;
wire slo__sro_n611;
wire slo__sro_n612;
wire slo__sro_n613;
wire slo__sro_n727;
wire slo__sro_n728;
wire slo__sro_n490;
wire slo__sro_n491;
wire slo__sro_n492;
wire slo__sro_n493;
wire slo__sro_n729;
wire slo__sro_n730;
wire opt_ipo_n1278;
wire CLOCK_slo__sro_n1332;
wire CLOCK_slo__sro_n1333;
wire CLOCK_slo__sro_n1334;
wire CLOCK_slo__mro_n1354;
wire CLOCK_slo__sro_n1383;
wire CLOCK_slo__sro_n1384;
wire CLOCK_slo__mro_n1394;
wire CLOCK_slo__sro_n1432;
wire CLOCK_slo__sro_n1433;
wire CLOCK_slo__sro_n1434;
wire CLOCK_slo__sro_n1435;
wire CLOCK_slo__sro_n1465;
wire CLOCK_slo__sro_n1466;
wire CLOCK_slo__sro_n1467;
wire CLOCK_slo__sro_n1468;
wire CLOCK_slo__xsl_n1522;
wire CLOCK_slo__xsl_n1523;
wire CLOCK_slo__sro_n1706;
wire CLOCK_slo__sro_n1769;
wire CLOCK_slo__sro_n1770;
wire CLOCK_slo__sro_n1771;
wire CLOCK_slo__sro_n1772;


INV_X1 i_36 (.ZN (n_34), .A (p_0[30]));
INV_X1 i_35 (.ZN (n_33), .A (p_1[30]));
INV_X2 i_34 (.ZN (n_32), .A (n_30));
INV_X1 slo__sro_c260 (.ZN (slo__sro_n366), .A (n_21));
NAND2_X1 CLOCK_slo__sro_c1189 (.ZN (CLOCK_slo__sro_n1771), .A1 (p_1[27]), .A2 (p_0[27]));
OAI22_X1 i_31 (.ZN (n_0), .A1 (n_34), .A2 (p_1[30]), .B1 (p_0[30]), .B2 (n_33));
XNOR2_X1 i_0 (.ZN (p_2[30]), .A (n_32), .B (n_0));
FA_X1 i_30 (.CO (n_30), .S (p_2[29]), .A (p_0[29]), .B (p_1[29]), .CI (n_29));
FA_X1 i_29 (.CO (n_29), .S (p_2[28]), .A (p_0[28]), .B (p_1[28]), .CI (CLOCK_slo__sro_n1769));
INV_X1 slo__sro_c45 (.ZN (slo__sro_n115), .A (n_15));
FA_X1 i_26 (.CO (n_26), .S (p_2[25]), .A (p_0[25]), .B (p_1[25]), .CI (n_25));
FA_X1 i_25 (.CO (n_25), .S (p_2[24]), .A (p_0[24]), .B (p_1[24]), .CI (CLOCK_slo__sro_n1466));
OAI21_X2 CLOCK_slo__sro_c1004 (.ZN (slo__n265), .A (slo__sro_n173), .B1 (slo__sro_n172), .B2 (slo__sro_n174));
INV_X1 slo__sro_c156 (.ZN (slo__sro_n225), .A (p_0[7]));
NAND2_X1 slo__sro_c311 (.ZN (slo__sro_n441), .A1 (p_1[17]), .A2 (p_0[17]));
XNOR2_X2 CLOCK_slo__mro_c857 (.ZN (CLOCK_slo__mro_n1394), .A (p_1[22]), .B (p_0[22]));
FA_X1 i_20 (.CO (n_20), .S (p_2[19]), .A (p_0[19]), .B (p_1[19]), .CI (n_19));
OAI21_X1 slo__sro_c489 (.ZN (n_6), .A (slo__sro_n729), .B1 (slo__sro_n730), .B2 (slo__sro_n728));
NOR2_X1 slo__sro_c429 (.ZN (slo__sro_n611), .A1 (p_1[10]), .A2 (p_0[10]));
INV_X1 slo__sro_c29 (.ZN (slo__sro_n97), .A (n_26));
INV_X1 slo__sro_c76 (.ZN (slo__sro_n146), .A (slo__sro_n363));
INV_X1 CLOCK_slo__sro_c843 (.ZN (CLOCK_slo__sro_n1384), .A (n_20));
FA_X1 i_14 (.CO (n_14), .S (p_2[13]), .A (p_0[13]), .B (p_1[13]), .CI (n_13));
INV_X1 slo__sro_c15 (.ZN (slo__sro_n80), .A (n_16));
NAND2_X1 slo__sro_c261 (.ZN (slo__sro_n365), .A1 (p_1[21]), .A2 (p_0[21]));
INV_X1 slo__sro_c486 (.ZN (slo__sro_n730), .A (n_5));
FA_X1 i_10 (.CO (n_10), .S (p_2[9]), .A (p_0[9]), .B (p_1[9]), .CI (n_9));
FA_X1 i_9 (.CO (n_9), .S (p_2[8]), .A (p_0[8]), .B (p_1[8]), .CI (opt_ipo_n1278));
INV_X1 slo__sro_c172 (.ZN (slo__sro_n241), .A (n_30));
XNOR2_X1 slo__sro_c162 (.ZN (p_2[7]), .A (slo__sro_n220), .B (p_1[7]));
XNOR2_X1 CLOCK_slo__mro_c779 (.ZN (CLOCK_slo__mro_n1314), .A (p_1[17]), .B (p_0[17]));
FA_X1 i_5 (.CO (n_5), .S (p_2[4]), .A (p_0[4]), .B (p_1[4]), .CI (n_4));
FA_X1 i_4 (.CO (n_4), .S (p_2[3]), .A (p_0[3]), .B (p_1[3]), .CI (CLOCK_slo__sro_n1432));
FA_X1 i_2 (.CO (n_2), .S (p_2[1]), .A (p_0[1]), .B (p_1[1]), .CI (n_1));
HA_X1 i_1 (.CO (n_1), .S (p_2[0]), .A (p_0[0]), .B (p_1[0]));
INV_X1 slo__sro_c1 (.ZN (slo__sro_n66), .A (n_12));
NAND2_X1 slo__sro_c2 (.ZN (slo__sro_n65), .A1 (p_1[12]), .A2 (p_0[12]));
NOR2_X1 slo__sro_c3 (.ZN (slo__sro_n64), .A1 (p_1[12]), .A2 (p_0[12]));
OAI21_X1 slo__sro_c4 (.ZN (n_13), .A (slo__sro_n65), .B1 (slo__sro_n66), .B2 (slo__sro_n64));
XNOR2_X1 slo__sro_c5 (.ZN (slo__sro_n63), .A (p_1[12]), .B (p_0[12]));
XNOR2_X1 slo__sro_c6 (.ZN (p_2[12]), .A (slo__sro_n63), .B (n_12));
NAND2_X1 slo__sro_c16 (.ZN (slo__sro_n79), .A1 (p_1[16]), .A2 (p_0[16]));
NOR2_X1 slo__sro_c17 (.ZN (slo__sro_n78), .A1 (p_1[16]), .A2 (p_0[16]));
OAI21_X2 slo__sro_c18 (.ZN (slo__sro_n77), .A (slo__sro_n79), .B1 (slo__sro_n80), .B2 (slo__sro_n78));
XNOR2_X1 slo__sro_c19 (.ZN (slo__sro_n76), .A (p_1[16]), .B (p_0[16]));
XNOR2_X2 slo__sro_c20 (.ZN (p_2[16]), .A (slo__sro_n76), .B (CLOCK_slo__xsl_n1522));
NAND2_X1 slo__sro_c30 (.ZN (slo__sro_n96), .A1 (p_1[26]), .A2 (p_0[26]));
NOR2_X1 slo__sro_c31 (.ZN (slo__sro_n95), .A1 (p_1[26]), .A2 (p_0[26]));
OAI21_X1 slo__sro_c32 (.ZN (slo__sro_n94), .A (slo__sro_n96), .B1 (slo__sro_n97), .B2 (slo__sro_n95));
XNOR2_X1 slo__sro_c33 (.ZN (slo__sro_n93), .A (p_1[26]), .B (p_0[26]));
XNOR2_X1 slo__sro_c34 (.ZN (p_2[26]), .A (slo__sro_n93), .B (n_26));
NAND2_X1 slo__sro_c46 (.ZN (slo__sro_n114), .A1 (p_1[15]), .A2 (p_0[15]));
NOR2_X2 slo__sro_c47 (.ZN (slo__sro_n113), .A1 (p_1[15]), .A2 (p_0[15]));
OAI21_X2 slo__sro_c48 (.ZN (n_16), .A (slo__sro_n114), .B1 (slo__sro_n115), .B2 (slo__sro_n113));
XNOR2_X2 slo__sro_c49 (.ZN (slo__sro_n112), .A (p_1[15]), .B (p_0[15]));
XNOR2_X1 slo__sro_c50 (.ZN (p_2[15]), .A (slo__sro_n112), .B (n_15));
OAI21_X1 CLOCK_slo__sro_c846 (.ZN (n_21), .A (CLOCK_slo__sro_n1383), .B1 (CLOCK_slo__sro_n1384), .B2 (CLOCK_slo__sro_n1382));
NOR2_X1 slo__sro_c78 (.ZN (slo__sro_n144), .A1 (p_1[22]), .A2 (p_0[22]));
OAI21_X1 slo__sro_c79 (.ZN (slo__sro_n143), .A (CLOCK_slo__mro_n1354), .B1 (slo__sro_n146), .B2 (slo__sro_n144));
INV_X1 CLOCK_slo__sro_c898 (.ZN (CLOCK_slo__sro_n1435), .A (n_2));
NAND2_X1 CLOCK_slo__sro_c899 (.ZN (CLOCK_slo__sro_n1434), .A1 (p_1[2]), .A2 (p_0[2]));
INV_X2 slo__sro_c157 (.ZN (slo__sro_n224), .A (slo__n265));
NAND2_X2 slo__sro_c158 (.ZN (slo__sro_n223), .A1 (slo__sro_n224), .A2 (slo__sro_n225));
AOI22_X4 slo__sro_c159 (.ZN (slo__sro_n222), .A1 (slo__sro_n223), .A2 (p_1[7]), .B1 (n_7), .B2 (p_0[7]));
XNOR2_X1 CLOCK_slo__mro_c780 (.ZN (p_2[17]), .A (CLOCK_slo__mro_n1314), .B (slo__sro_n77));
XNOR2_X1 slo__sro_c161 (.ZN (slo__sro_n220), .A (n_7), .B (p_0[7]));
INV_X1 slo__sro_c103 (.ZN (slo__sro_n174), .A (n_6));
NAND2_X1 slo__sro_c104 (.ZN (slo__sro_n173), .A1 (p_1[6]), .A2 (p_0[6]));
NOR2_X2 slo__sro_c105 (.ZN (slo__sro_n172), .A1 (p_1[6]), .A2 (p_0[6]));
OAI21_X2 slo__sro_c106 (.ZN (n_7), .A (slo__sro_n173), .B1 (slo__sro_n174), .B2 (slo__sro_n172));
XNOR2_X2 slo__sro_c107 (.ZN (slo__sro_n171), .A (p_1[6]), .B (p_0[6]));
XNOR2_X2 slo__sro_c108 (.ZN (p_2[6]), .A (slo__sro_n171), .B (n_6));
NOR2_X1 slo__sro_c173 (.ZN (slo__sro_n240), .A1 (n_33), .A2 (p_0[30]));
NAND2_X1 slo__sro_c174 (.ZN (slo__sro_n239), .A1 (slo__sro_n240), .A2 (slo__sro_n241));
OR2_X1 slo__sro_c175 (.ZN (slo__sro_n238), .A1 (p_1[30]), .A2 (n_34));
OAI21_X1 slo__sro_c176 (.ZN (slo__sro_n237), .A (slo__sro_n239), .B1 (n_32), .B2 (slo__sro_n238));
INV_X1 slo__sro_c232 (.ZN (slo__sro_n312), .A (slo__sro_n610));
INV_X1 slo__sro_c310 (.ZN (slo__sro_n442), .A (slo__sro_n77));
INV_X1 CLOCK_slo__sro_c1188 (.ZN (CLOCK_slo__sro_n1772), .A (slo__sro_n94));
NAND2_X1 slo__sro_c428 (.ZN (slo__sro_n612), .A1 (p_1[10]), .A2 (p_0[10]));
INV_X2 slo__sro_c427 (.ZN (slo__sro_n613), .A (n_10));
NAND2_X1 slo__sro_c233 (.ZN (slo__sro_n311), .A1 (p_1[11]), .A2 (p_0[11]));
NOR2_X1 slo__sro_c234 (.ZN (slo__sro_n310), .A1 (p_1[11]), .A2 (p_0[11]));
OAI21_X2 slo__sro_c235 (.ZN (n_12), .A (slo__sro_n311), .B1 (slo__sro_n312), .B2 (slo__sro_n310));
XNOR2_X1 slo__sro_c236 (.ZN (slo__sro_n309), .A (p_1[11]), .B (p_0[11]));
XNOR2_X1 slo__sro_c237 (.ZN (p_2[11]), .A (slo__sro_n610), .B (slo__sro_n309));
NOR2_X1 slo__sro_c262 (.ZN (slo__sro_n364), .A1 (p_1[21]), .A2 (p_0[21]));
OAI21_X1 slo__sro_c263 (.ZN (slo__sro_n363), .A (slo__sro_n365), .B1 (slo__sro_n366), .B2 (slo__sro_n364));
XNOR2_X1 slo__sro_c264 (.ZN (slo__sro_n362), .A (p_1[21]), .B (p_0[21]));
XNOR2_X1 slo__sro_c265 (.ZN (p_2[21]), .A (n_21), .B (slo__sro_n362));
NOR2_X1 slo__sro_c312 (.ZN (slo__sro_n440), .A1 (p_1[17]), .A2 (p_0[17]));
OAI21_X2 slo__sro_c313 (.ZN (slo__sro_n439), .A (slo__sro_n441), .B1 (slo__sro_n440), .B2 (slo__sro_n442));
INV_X1 CLOCK_slo__sro_c793 (.ZN (CLOCK_slo__sro_n1334), .A (n_14));
NAND2_X1 CLOCK_slo__sro_c794 (.ZN (CLOCK_slo__sro_n1333), .A1 (p_1[14]), .A2 (p_0[14]));
OAI21_X2 slo__sro_c430 (.ZN (slo__sro_n610), .A (slo__sro_n612), .B1 (slo__sro_n613), .B2 (slo__sro_n611));
XNOR2_X1 slo__sro_c431 (.ZN (slo__sro_n609), .A (p_1[10]), .B (p_0[10]));
XNOR2_X1 slo__sro_c432 (.ZN (p_2[10]), .A (n_10), .B (slo__sro_n609));
NAND2_X1 slo__sro_c487 (.ZN (slo__sro_n729), .A1 (p_1[5]), .A2 (p_0[5]));
NOR2_X1 slo__sro_c488 (.ZN (slo__sro_n728), .A1 (p_1[5]), .A2 (p_0[5]));
INV_X1 slo__sro_c366 (.ZN (slo__sro_n493), .A (slo__sro_n439));
NAND2_X1 slo__sro_c367 (.ZN (slo__sro_n492), .A1 (p_1[18]), .A2 (p_0[18]));
NOR2_X2 slo__sro_c368 (.ZN (slo__sro_n491), .A1 (p_1[18]), .A2 (p_0[18]));
OAI21_X2 slo__sro_c369 (.ZN (n_19), .A (slo__sro_n492), .B1 (slo__sro_n493), .B2 (slo__sro_n491));
XNOR2_X1 slo__sro_c370 (.ZN (slo__sro_n490), .A (p_1[18]), .B (p_0[18]));
XNOR2_X1 slo__sro_c371 (.ZN (p_2[18]), .A (slo__sro_n490), .B (slo__sro_n439));
XNOR2_X1 slo__sro_c490 (.ZN (slo__sro_n727), .A (p_1[5]), .B (p_0[5]));
XNOR2_X1 slo__sro_c491 (.ZN (p_2[5]), .A (n_5), .B (slo__sro_n727));
NOR2_X1 CLOCK_slo__sro_c845 (.ZN (CLOCK_slo__sro_n1382), .A1 (p_1[20]), .A2 (p_0[20]));
INV_X2 opt_ipo_c750 (.ZN (opt_ipo_n1278), .A (slo__sro_n222));
NOR2_X1 CLOCK_slo__sro_c795 (.ZN (CLOCK_slo__sro_n1332), .A1 (p_1[14]), .A2 (p_0[14]));
OAI21_X2 CLOCK_slo__sro_c796 (.ZN (n_15), .A (CLOCK_slo__sro_n1333), .B1 (CLOCK_slo__sro_n1334), .B2 (CLOCK_slo__sro_n1332));
XNOR2_X1 CLOCK_slo__sro_c797 (.ZN (CLOCK_slo__sro_n1331), .A (p_1[14]), .B (p_0[14]));
XNOR2_X1 CLOCK_slo__sro_c798 (.ZN (p_2[14]), .A (n_14), .B (CLOCK_slo__sro_n1331));
NAND2_X1 CLOCK_slo__sro_c844 (.ZN (CLOCK_slo__sro_n1383), .A1 (p_1[20]), .A2 (p_0[20]));
NAND2_X1 CLOCK_slo__mro_c818 (.ZN (CLOCK_slo__mro_n1354), .A1 (p_1_22_PP_5), .A2 (p_0[22]));
XNOR2_X1 CLOCK_slo__sro_c847 (.ZN (CLOCK_slo__sro_n1381), .A (p_1[20]), .B (p_0[20]));
XNOR2_X1 CLOCK_slo__sro_c848 (.ZN (p_2[20]), .A (CLOCK_slo__sro_n1381), .B (n_20));
XNOR2_X2 CLOCK_slo__mro_c858 (.ZN (p_2[22]), .A (CLOCK_slo__mro_n1394), .B (slo__sro_n363));
NOR2_X1 CLOCK_slo__sro_c900 (.ZN (CLOCK_slo__sro_n1433), .A1 (p_1[2]), .A2 (p_0[2]));
OAI21_X1 CLOCK_slo__sro_c901 (.ZN (CLOCK_slo__sro_n1432), .A (CLOCK_slo__sro_n1434)
    , .B1 (CLOCK_slo__sro_n1435), .B2 (CLOCK_slo__sro_n1433));
XNOR2_X1 CLOCK_slo__sro_c902 (.ZN (CLOCK_slo__sro_n1431), .A (p_1[2]), .B (p_0[2]));
XNOR2_X1 CLOCK_slo__sro_c903 (.ZN (p_2[2]), .A (n_2), .B (CLOCK_slo__sro_n1431));
NAND2_X1 CLOCK_slo__sro_c928 (.ZN (CLOCK_slo__sro_n1468), .A1 (slo__sro_n143), .A2 (p_0[23]));
OAI21_X1 CLOCK_slo__sro_c929 (.ZN (CLOCK_slo__sro_n1467), .A (p_1[23]), .B1 (slo__sro_n143), .B2 (p_0[23]));
NAND2_X1 CLOCK_slo__sro_c930 (.ZN (CLOCK_slo__sro_n1466), .A1 (CLOCK_slo__sro_n1468), .A2 (CLOCK_slo__sro_n1467));
XNOR2_X1 CLOCK_slo__sro_c931 (.ZN (CLOCK_slo__sro_n1465), .A (p_1[23]), .B (p_0[23]));
XNOR2_X1 CLOCK_slo__sro_c932 (.ZN (p_2[23]), .A (CLOCK_slo__sro_n1465), .B (slo__sro_n143));
INV_X1 CLOCK_slo__sro_c1126 (.ZN (CLOCK_slo__sro_n1706), .A (p_0[31]));
INV_X1 CLOCK_slo__xsl_c974 (.ZN (CLOCK_slo__xsl_n1523), .A (n_16));
INV_X1 CLOCK_slo__xsl_c975 (.ZN (CLOCK_slo__xsl_n1522), .A (CLOCK_slo__xsl_n1523));
XNOR2_X1 CLOCK_slo__sro_c1127 (.ZN (p_2[31]), .A (slo__sro_n237), .B (CLOCK_slo__sro_n1706));
NOR2_X1 CLOCK_slo__sro_c1190 (.ZN (CLOCK_slo__sro_n1770), .A1 (p_1[27]), .A2 (p_0[27]));
OAI21_X1 CLOCK_slo__sro_c1191 (.ZN (CLOCK_slo__sro_n1769), .A (CLOCK_slo__sro_n1771)
    , .B1 (CLOCK_slo__sro_n1772), .B2 (CLOCK_slo__sro_n1770));
XNOR2_X1 CLOCK_slo__sro_c1192 (.ZN (CLOCK_slo__sro_n1768), .A (p_1[27]), .B (p_0[27]));
XNOR2_X1 CLOCK_slo__sro_c1193 (.ZN (p_2[27]), .A (CLOCK_slo__sro_n1768), .B (slo__sro_n94));

endmodule //datapath__0_227

module datapath__0_226 (p_0_24_PP_1, Multiplier, p_0, p_1);

output [31:0] p_1;
input [31:0] Multiplier;
input [31:0] p_0;
input p_0_24_PP_1;
wire CLOCK_slo__sro_n1549;
wire slo__sro_n604;
wire n_1;
wire n_2;
wire n_3;
wire n_4;
wire n_5;
wire n_6;
wire n_7;
wire n_8;
wire n_9;
wire n_10;
wire n_11;
wire n_14;
wire n_15;
wire n_16;
wire slo__sro_n297;
wire slo__sro_n462;
wire n_20;
wire n_23;
wire n_25;
wire n_27;
wire n_28;
wire n_29;
wire n_30;
wire n_32;
wire n_0;
wire n_34;
wire n_33;
wire slo__sro_n59;
wire slo__sro_n60;
wire slo__sro_n61;
wire slo__sro_n62;
wire slo__sro_n63;
wire slo__sro_n76;
wire slo__sro_n78;
wire slo__sro_n79;
wire slo__sro_n80;
wire slo__sro_n93;
wire slo__sro_n94;
wire slo__sro_n95;
wire slo__sro_n96;
wire slo__sro_n97;
wire slo__sro_n110;
wire slo__sro_n111;
wire slo__sro_n112;
wire slo__sro_n113;
wire slo__sro_n155;
wire slo__sro_n156;
wire slo__sro_n157;
wire slo__sro_n158;
wire slo__sro_n159;
wire slo__sro_n174;
wire slo__sro_n175;
wire slo__sro_n176;
wire slo__sro_n177;
wire slo__sro_n178;
wire slo__sro_n253;
wire slo__sro_n254;
wire slo__sro_n255;
wire slo__sro_n256;
wire slo__sro_n266;
wire slo__sro_n267;
wire slo__sro_n268;
wire slo__sro_n269;
wire slo__sro_n279;
wire slo__sro_n280;
wire slo__sro_n281;
wire slo__sro_n282;
wire slo__sro_n294;
wire slo__sro_n295;
wire slo__sro_n296;
wire slo__sro_n236;
wire slo__sro_n237;
wire slo__sro_n238;
wire slo__sro_n239;
wire slo__sro_n240;
wire slo__sro_n298;
wire slo__sro_n570;
wire slo__sro_n810;
wire slo__sro_n571;
wire slo__sro_n572;
wire slo__sro_n573;
wire slo__sro_n574;
wire slo__sro_n605;
wire slo__sro_n606;
wire slo__sro_n622;
wire slo__sro_n623;
wire slo__sro_n624;
wire slo__sro_n811;
wire slo__sro_n812;
wire CLOCK_slo__mro_n1532;
wire slo__n878;
wire slo__sro_n907;
wire slo__sro_n908;
wire slo__sro_n909;
wire slo__sro_n910;
wire CLOCK_slo__sro_n1550;
wire CLOCK_slo__sro_n1551;
wire CLOCK_slo__sro_n1552;
wire CLOCK_slo__sro_n1562;
wire CLOCK_slo__sro_n1563;
wire CLOCK_slo__sro_n1564;
wire CLOCK_slo__sro_n1565;
wire CLOCK_slo__sro_n1566;
wire CLOCK_slo__sro_n1653;
wire CLOCK_slo__sro_n1654;
wire CLOCK_slo__sro_n1655;
wire CLOCK_slo__sro_n1656;
wire CLOCK_slo__sro_n1668;
wire CLOCK_slo__sro_n1669;
wire CLOCK_slo__sro_n1670;
wire CLOCK_slo__sro_n1671;
wire CLOCK_slo__sro_n2036;
wire CLOCK_slo__sro_n2037;
wire CLOCK_slo__sro_n2038;
wire CLOCK_slo__sro_n2039;
wire CLOCK_slo__sro_n2040;


INV_X1 i_36 (.ZN (n_34), .A (Multiplier[30]));
INV_X1 i_35 (.ZN (n_33), .A (p_0[30]));
INV_X2 i_34 (.ZN (n_32), .A (n_30));
XOR2_X1 i_32 (.Z (p_1[31]), .A (CLOCK_slo__sro_n1562), .B (Multiplier[31]));
OAI22_X1 i_31 (.ZN (n_0), .A1 (n_34), .A2 (p_0[30]), .B1 (n_33), .B2 (Multiplier[30]));
XNOR2_X1 i_0 (.ZN (p_1[30]), .A (n_32), .B (n_0));
FA_X1 i_30 (.CO (n_30), .S (p_1[29]), .A (Multiplier[29]), .B (p_0[29]), .CI (n_29));
INV_X1 slo__sro_c208 (.ZN (slo__sro_n298), .A (slo__sro_n237));
XNOR2_X2 CLOCK_slo__mro_c1019 (.ZN (p_1[6]), .A (CLOCK_slo__mro_n1532), .B (n_6));
INV_X2 slo__sro_c83 (.ZN (slo__sro_n159), .A (n_23));
INV_X1 slo__sro_c15 (.ZN (slo__sro_n80), .A (n_20));
INV_X1 slo__sro_c425 (.ZN (slo__sro_n624), .A (p_0[6]));
INV_X1 slo__sro_c99 (.ZN (slo__sro_n178), .A (n_11));
FA_X1 i_23 (.CO (n_23), .S (p_1[22]), .A (Multiplier[22]), .B (p_0[22]), .CI (slo__sro_n571));
NAND2_X1 slo__sro_c410 (.ZN (slo__sro_n606), .A1 (slo__sro_n156), .A2 (Multiplier[24]));
INV_X1 slo__sro_c29 (.ZN (slo__sro_n97), .A (slo__sro_n175));
FA_X1 i_20 (.CO (n_20), .S (p_1[19]), .A (Multiplier[19]), .B (p_0[19]), .CI (CLOCK_slo__sro_n2037));
OAI21_X2 slo__sro_c320 (.ZN (slo__sro_n462), .A (slo__sro_n79), .B1 (slo__sro_n80), .B2 (slo__sro_n78));
OAI21_X2 slo__sro_c211 (.ZN (slo__sro_n295), .A (slo__sro_n297), .B1 (slo__sro_n298), .B2 (slo__sro_n296));
NOR2_X1 CLOCK_slo__sro_c1034 (.ZN (CLOCK_slo__sro_n1550), .A1 (n_1), .A2 (Multiplier[1]));
FA_X1 i_15 (.CO (n_15), .S (p_1[14]), .A (Multiplier[14]), .B (p_0[14]), .CI (n_14));
FA_X1 i_14 (.CO (n_14), .S (p_1[13]), .A (Multiplier[13]), .B (p_0[13]), .CI (slo__sro_n94));
INV_X1 slo__sro_c43 (.ZN (slo__sro_n113), .A (p_0[26]));
INV_X1 slo__sro_c166 (.ZN (slo__sro_n256), .A (n_2));
INV_X1 CLOCK_slo__sro_c1503 (.ZN (CLOCK_slo__sro_n2040), .A (slo__sro_n295));
FA_X1 i_10 (.CO (n_10), .S (p_1[9]), .A (Multiplier[9]), .B (p_0[9]), .CI (n_9));
FA_X1 i_9 (.CO (n_9), .S (p_1[8]), .A (Multiplier[8]), .B (p_0[8]), .CI (n_8));
INV_X1 slo__sro_c194 (.ZN (slo__sro_n282), .A (n_28));
NAND2_X1 slo__sro_c566 (.ZN (n_28), .A1 (slo__sro_n811), .A2 (slo__sro_n812));
INV_X1 CLOCK_slo__sro_c1172 (.ZN (CLOCK_slo__sro_n1671), .A (n_10));
FA_X1 i_5 (.CO (n_5), .S (p_1[4]), .A (Multiplier[4]), .B (p_0[4]), .CI (n_4));
FA_X1 i_4 (.CO (n_4), .S (p_1[3]), .A (Multiplier[3]), .B (p_0[3]), .CI (n_3));
INV_X1 slo__sro_c180 (.ZN (slo__sro_n269), .A (n_7));
INV_X1 CLOCK_slo__sro_c1048 (.ZN (CLOCK_slo__sro_n1566), .A (n_30));
HA_X1 i_1 (.CO (n_1), .S (p_1[0]), .A (Multiplier[0]), .B (p_0[0]));
INV_X1 slo__sro_c1 (.ZN (slo__sro_n63), .A (n_25));
NAND2_X1 slo__sro_c2 (.ZN (slo__sro_n62), .A1 (p_0[25]), .A2 (Multiplier[25]));
NOR2_X2 slo__sro_c3 (.ZN (slo__sro_n61), .A1 (p_0[25]), .A2 (Multiplier[25]));
OAI21_X2 slo__sro_c4 (.ZN (slo__sro_n60), .A (slo__sro_n62), .B1 (slo__sro_n61), .B2 (slo__sro_n63));
XNOR2_X2 slo__sro_c5 (.ZN (slo__sro_n59), .A (p_0[25]), .B (Multiplier[25]));
XNOR2_X1 slo__sro_c6 (.ZN (p_1[25]), .A (slo__sro_n59), .B (n_25));
NAND2_X1 slo__sro_c16 (.ZN (slo__sro_n79), .A1 (p_0[20]), .A2 (Multiplier[20]));
NOR2_X1 slo__sro_c17 (.ZN (slo__sro_n78), .A1 (p_0[20]), .A2 (Multiplier[20]));
INV_X1 slo__sro_c635 (.ZN (slo__sro_n910), .A (n_15));
XNOR2_X2 slo__sro_c19 (.ZN (slo__sro_n76), .A (p_0[20]), .B (Multiplier[20]));
XNOR2_X1 slo__sro_c20 (.ZN (p_1[20]), .A (n_20), .B (slo__sro_n76));
NAND2_X1 slo__sro_c30 (.ZN (slo__sro_n96), .A1 (p_0[12]), .A2 (Multiplier[12]));
NOR2_X1 slo__sro_c31 (.ZN (slo__sro_n95), .A1 (p_0[12]), .A2 (Multiplier[12]));
OAI21_X1 slo__sro_c32 (.ZN (slo__sro_n94), .A (slo__sro_n96), .B1 (slo__sro_n97), .B2 (slo__sro_n95));
XNOR2_X1 slo__sro_c33 (.ZN (slo__sro_n93), .A (p_0[12]), .B (Multiplier[12]));
XNOR2_X1 slo__sro_c34 (.ZN (p_1[12]), .A (slo__sro_n93), .B (slo__sro_n175));
NAND2_X1 slo__sro_c44 (.ZN (slo__sro_n112), .A1 (slo__sro_n60), .A2 (Multiplier[26]));
NOR2_X1 slo__sro_c45 (.ZN (slo__sro_n111), .A1 (slo__sro_n60), .A2 (Multiplier[26]));
OAI21_X2 slo__sro_c46 (.ZN (n_27), .A (slo__sro_n112), .B1 (slo__sro_n113), .B2 (slo__sro_n111));
XNOR2_X2 slo__sro_c47 (.ZN (slo__sro_n110), .A (slo__sro_n60), .B (Multiplier[26]));
XNOR2_X2 slo__sro_c48 (.ZN (p_1[26]), .A (slo__sro_n110), .B (p_0[26]));
NAND2_X1 slo__sro_c84 (.ZN (slo__sro_n158), .A1 (p_0[23]), .A2 (Multiplier[23]));
NOR2_X1 slo__sro_c85 (.ZN (slo__sro_n157), .A1 (p_0[23]), .A2 (Multiplier[23]));
OAI21_X2 slo__sro_c86 (.ZN (slo__sro_n156), .A (slo__sro_n158), .B1 (slo__sro_n159), .B2 (slo__sro_n157));
XNOR2_X2 slo__sro_c87 (.ZN (slo__sro_n155), .A (p_0[23]), .B (Multiplier[23]));
XNOR2_X1 slo__sro_c88 (.ZN (p_1[23]), .A (slo__sro_n155), .B (n_23));
NAND2_X1 slo__sro_c100 (.ZN (slo__sro_n177), .A1 (p_0[11]), .A2 (Multiplier[11]));
NOR2_X1 slo__sro_c101 (.ZN (slo__sro_n176), .A1 (p_0[11]), .A2 (Multiplier[11]));
OAI21_X2 slo__sro_c102 (.ZN (slo__sro_n175), .A (slo__sro_n177), .B1 (slo__sro_n176), .B2 (slo__sro_n178));
XNOR2_X1 slo__sro_c103 (.ZN (slo__sro_n174), .A (p_0[11]), .B (Multiplier[11]));
XNOR2_X1 slo__sro_c104 (.ZN (p_1[11]), .A (slo__sro_n174), .B (n_11));
NAND2_X1 slo__sro_c167 (.ZN (slo__sro_n255), .A1 (p_0[2]), .A2 (Multiplier[2]));
NOR2_X1 slo__sro_c168 (.ZN (slo__sro_n254), .A1 (p_0[2]), .A2 (Multiplier[2]));
OAI21_X1 slo__sro_c169 (.ZN (n_3), .A (slo__sro_n255), .B1 (slo__sro_n256), .B2 (slo__sro_n254));
XNOR2_X2 slo__sro_c170 (.ZN (slo__sro_n253), .A (p_0[2]), .B (Multiplier[2]));
XNOR2_X2 slo__sro_c171 (.ZN (p_1[2]), .A (slo__sro_n253), .B (n_2));
NAND2_X1 slo__sro_c181 (.ZN (slo__sro_n268), .A1 (p_0[7]), .A2 (Multiplier[7]));
NOR2_X1 slo__sro_c182 (.ZN (slo__sro_n267), .A1 (p_0[7]), .A2 (Multiplier[7]));
OAI21_X1 slo__sro_c183 (.ZN (n_8), .A (slo__sro_n268), .B1 (slo__sro_n267), .B2 (slo__sro_n269));
XNOR2_X1 slo__sro_c184 (.ZN (slo__sro_n266), .A (p_0[7]), .B (Multiplier[7]));
XNOR2_X1 slo__sro_c185 (.ZN (p_1[7]), .A (slo__sro_n266), .B (n_7));
NAND2_X1 slo__sro_c195 (.ZN (slo__sro_n281), .A1 (p_0[28]), .A2 (Multiplier[28]));
NOR2_X2 slo__sro_c196 (.ZN (slo__sro_n280), .A1 (p_0[28]), .A2 (Multiplier[28]));
OAI21_X1 slo__sro_c197 (.ZN (n_29), .A (slo__sro_n281), .B1 (slo__sro_n280), .B2 (slo__sro_n282));
XNOR2_X1 slo__sro_c198 (.ZN (slo__sro_n279), .A (p_0[28]), .B (Multiplier[28]));
XNOR2_X1 slo__sro_c199 (.ZN (p_1[28]), .A (slo__sro_n279), .B (n_28));
NAND2_X1 slo__sro_c209 (.ZN (slo__sro_n297), .A1 (p_0[17]), .A2 (Multiplier[17]));
NOR2_X1 slo__sro_c210 (.ZN (slo__sro_n296), .A1 (p_0[17]), .A2 (Multiplier[17]));
INV_X2 slo__sro_c152 (.ZN (slo__sro_n240), .A (n_16));
NAND2_X1 slo__sro_c153 (.ZN (slo__sro_n239), .A1 (p_0[16]), .A2 (Multiplier[16]));
NOR2_X2 slo__sro_c154 (.ZN (slo__sro_n238), .A1 (p_0[16]), .A2 (Multiplier[16]));
OAI21_X2 slo__sro_c155 (.ZN (slo__sro_n237), .A (slo__sro_n239), .B1 (slo__sro_n240), .B2 (slo__sro_n238));
XNOR2_X1 slo__sro_c156 (.ZN (slo__sro_n236), .A (p_0[16]), .B (Multiplier[16]));
XNOR2_X1 slo__sro_c157 (.ZN (p_1[16]), .A (n_16), .B (slo__sro_n236));
XNOR2_X2 slo__sro_c212 (.ZN (slo__sro_n294), .A (p_0[17]), .B (Multiplier[17]));
INV_X1 slo__sro_c387 (.ZN (slo__sro_n574), .A (slo__sro_n462));
NAND2_X1 slo__sro_c388 (.ZN (slo__sro_n573), .A1 (p_0[21]), .A2 (Multiplier[21]));
OAI21_X1 slo__sro_c565 (.ZN (slo__sro_n811), .A (p_0[27]), .B1 (n_27), .B2 (Multiplier[27]));
NAND2_X1 slo__sro_c564 (.ZN (slo__sro_n812), .A1 (n_27), .A2 (Multiplier[27]));
NOR2_X1 slo__sro_c389 (.ZN (slo__sro_n572), .A1 (p_0[21]), .A2 (Multiplier[21]));
OAI21_X2 slo__sro_c390 (.ZN (slo__sro_n571), .A (slo__sro_n573), .B1 (slo__sro_n574), .B2 (slo__sro_n572));
XNOR2_X1 slo__sro_c391 (.ZN (slo__sro_n570), .A (p_0[21]), .B (Multiplier[21]));
XNOR2_X1 slo__sro_c392 (.ZN (p_1[21]), .A (slo__sro_n570), .B (slo__sro_n462));
NOR2_X1 slo__sro_c411 (.ZN (slo__sro_n605), .A1 (slo__sro_n156), .A2 (Multiplier[24]));
OAI21_X1 slo__sro_c412 (.ZN (n_25), .A (slo__sro_n606), .B1 (slo__sro_n605), .B2 (slo__n878));
XNOR2_X2 slo__sro_c413 (.ZN (slo__sro_n604), .A (slo__sro_n156), .B (Multiplier[24]));
XNOR2_X2 slo__sro_c414 (.ZN (p_1[24]), .A (slo__sro_n604), .B (p_0[24]));
NAND2_X1 slo__sro_c426 (.ZN (slo__sro_n623), .A1 (n_6), .A2 (Multiplier[6]));
NOR2_X1 slo__sro_c427 (.ZN (slo__sro_n622), .A1 (n_6), .A2 (Multiplier[6]));
OAI21_X1 slo__sro_c428 (.ZN (n_7), .A (slo__sro_n623), .B1 (slo__sro_n624), .B2 (slo__sro_n622));
INV_X1 CLOCK_slo__sro_c1032 (.ZN (CLOCK_slo__sro_n1552), .A (p_0[1]));
NAND2_X1 CLOCK_slo__sro_c1033 (.ZN (CLOCK_slo__sro_n1551), .A1 (n_1), .A2 (Multiplier[1]));
XNOR2_X1 slo__sro_c567 (.ZN (slo__sro_n810), .A (n_27), .B (Multiplier[27]));
XNOR2_X1 slo__sro_c568 (.ZN (p_1[27]), .A (slo__sro_n810), .B (p_0[27]));
XNOR2_X2 CLOCK_slo__mro_c1018 (.ZN (CLOCK_slo__mro_n1532), .A (p_0[6]), .B (Multiplier[6]));
INV_X1 slo__L2_c3_c623 (.ZN (slo__n878), .A (p_0_24_PP_1));
NAND2_X1 slo__sro_c636 (.ZN (slo__sro_n909), .A1 (p_0[15]), .A2 (Multiplier[15]));
NOR2_X1 slo__sro_c637 (.ZN (slo__sro_n908), .A1 (p_0[15]), .A2 (Multiplier[15]));
OAI21_X2 slo__sro_c638 (.ZN (n_16), .A (slo__sro_n909), .B1 (slo__sro_n910), .B2 (slo__sro_n908));
XNOR2_X1 slo__sro_c639 (.ZN (slo__sro_n907), .A (p_0[15]), .B (Multiplier[15]));
XNOR2_X1 slo__sro_c640 (.ZN (p_1[15]), .A (slo__sro_n907), .B (n_15));
OAI21_X1 CLOCK_slo__sro_c1035 (.ZN (n_2), .A (CLOCK_slo__sro_n1551), .B1 (CLOCK_slo__sro_n1552), .B2 (CLOCK_slo__sro_n1550));
XNOR2_X1 CLOCK_slo__sro_c1036 (.ZN (CLOCK_slo__sro_n1549), .A (n_1), .B (Multiplier[1]));
XNOR2_X1 CLOCK_slo__sro_c1037 (.ZN (p_1[1]), .A (CLOCK_slo__sro_n1549), .B (p_0[1]));
NOR2_X1 CLOCK_slo__sro_c1049 (.ZN (CLOCK_slo__sro_n1565), .A1 (n_33), .A2 (Multiplier[30]));
NAND2_X1 CLOCK_slo__sro_c1050 (.ZN (CLOCK_slo__sro_n1564), .A1 (CLOCK_slo__sro_n1566), .A2 (CLOCK_slo__sro_n1565));
OR2_X1 CLOCK_slo__sro_c1051 (.ZN (CLOCK_slo__sro_n1563), .A1 (p_0[30]), .A2 (n_34));
OAI21_X1 CLOCK_slo__sro_c1052 (.ZN (CLOCK_slo__sro_n1562), .A (CLOCK_slo__sro_n1564)
    , .B1 (n_32), .B2 (CLOCK_slo__sro_n1563));
INV_X1 CLOCK_slo__sro_c1156 (.ZN (CLOCK_slo__sro_n1656), .A (n_5));
NAND2_X1 CLOCK_slo__sro_c1157 (.ZN (CLOCK_slo__sro_n1655), .A1 (p_0[5]), .A2 (Multiplier[5]));
NOR2_X1 CLOCK_slo__sro_c1158 (.ZN (CLOCK_slo__sro_n1654), .A1 (p_0[5]), .A2 (Multiplier[5]));
OAI21_X2 CLOCK_slo__sro_c1159 (.ZN (n_6), .A (CLOCK_slo__sro_n1655), .B1 (CLOCK_slo__sro_n1654), .B2 (CLOCK_slo__sro_n1656));
XNOR2_X1 CLOCK_slo__sro_c1160 (.ZN (CLOCK_slo__sro_n1653), .A (p_0[5]), .B (Multiplier[5]));
XNOR2_X1 CLOCK_slo__sro_c1161 (.ZN (p_1[5]), .A (CLOCK_slo__sro_n1653), .B (n_5));
NAND2_X1 CLOCK_slo__sro_c1173 (.ZN (CLOCK_slo__sro_n1670), .A1 (p_0[10]), .A2 (Multiplier[10]));
NOR2_X1 CLOCK_slo__sro_c1174 (.ZN (CLOCK_slo__sro_n1669), .A1 (p_0[10]), .A2 (Multiplier[10]));
OAI21_X2 CLOCK_slo__sro_c1175 (.ZN (n_11), .A (CLOCK_slo__sro_n1670), .B1 (CLOCK_slo__sro_n1671), .B2 (CLOCK_slo__sro_n1669));
XNOR2_X1 CLOCK_slo__sro_c1176 (.ZN (CLOCK_slo__sro_n1668), .A (p_0[10]), .B (Multiplier[10]));
XNOR2_X1 CLOCK_slo__sro_c1177 (.ZN (p_1[10]), .A (CLOCK_slo__sro_n1668), .B (n_10));
XNOR2_X2 CLOCK_slo__mro_c1586 (.ZN (p_1[17]), .A (slo__sro_n294), .B (slo__sro_n237));
NAND2_X1 CLOCK_slo__sro_c1504 (.ZN (CLOCK_slo__sro_n2039), .A1 (p_0[18]), .A2 (Multiplier[18]));
NOR2_X1 CLOCK_slo__sro_c1505 (.ZN (CLOCK_slo__sro_n2038), .A1 (p_0[18]), .A2 (Multiplier[18]));
OAI21_X1 CLOCK_slo__sro_c1506 (.ZN (CLOCK_slo__sro_n2037), .A (CLOCK_slo__sro_n2039)
    , .B1 (CLOCK_slo__sro_n2040), .B2 (CLOCK_slo__sro_n2038));
XNOR2_X1 CLOCK_slo__sro_c1507 (.ZN (CLOCK_slo__sro_n2036), .A (p_0[18]), .B (Multiplier[18]));
XNOR2_X1 CLOCK_slo__sro_c1508 (.ZN (p_1[18]), .A (CLOCK_slo__sro_n2036), .B (slo__sro_n295));

endmodule //datapath__0_226

module datapath__0_222 (opt_ipoPP_5, p_0, p_1, p_2);

output [31:0] p_2;
input [31:0] p_0;
input [31:0] p_1;
input opt_ipoPP_5;
wire slo__sro_n558;
wire n_1;
wire n_2;
wire n_3;
wire n_4;
wire n_5;
wire n_6;
wire n_7;
wire n_8;
wire n_9;
wire n_10;
wire n_11;
wire n_12;
wire n_13;
wire n_14;
wire n_15;
wire n_16;
wire slo__sro_n932;
wire slo__sro_n195;
wire slo__sro_n698;
wire n_20;
wire n_21;
wire n_24;
wire n_25;
wire slo__sro_n433;
wire n_27;
wire n_28;
wire CLOCK_slo__sro_n1603;
wire n_30;
wire n_32;
wire n_0;
wire n_34;
wire n_33;
wire slo__sro_n180;
wire slo__sro_n181;
wire slo__sro_n182;
wire slo__sro_n183;
wire slo__sro_n80;
wire slo__sro_n81;
wire slo__sro_n82;
wire slo__sro_n83;
wire slo__sro_n84;
wire CLOCK_slo__xsl_n1812;
wire slo__sro_n197;
wire slo__sro_n198;
wire slo__sro_n199;
wire slo__sro_n933;
wire slo__sro_n557;
wire slo__sro_n429;
wire slo__sro_n430;
wire slo__sro_n431;
wire slo__sro_n333;
wire slo__sro_n334;
wire slo__sro_n335;
wire slo__sro_n336;
wire slo__sro_n432;
wire slo__sro_n374;
wire slo__sro_n375;
wire slo__sro_n376;
wire slo__sro_n377;
wire slo__sro_n378;
wire slo__sro_n559;
wire slo__sro_n560;
wire slo__sro_n561;
wire slo__sro_n697;
wire slo__sro_n530;
wire slo__sro_n531;
wire slo__sro_n532;
wire slo__sro_n533;
wire slo__sro_n534;
wire slo__sro_n699;
wire slo__sro_n700;
wire slo__sro_n934;
wire slo__sro_n915;
wire slo__sro_n916;
wire slo__sro_n917;
wire slo__sro_n918;
wire slo__sro_n962;
wire slo__sro_n963;
wire slo__sro_n964;
wire slo__sro_n965;
wire slo__sro_n975;
wire slo__sro_n976;
wire slo__sro_n977;
wire slo__sro_n978;
wire CLOCK_slo__sro_n1436;
wire CLOCK_slo__sro_n1437;
wire CLOCK_slo__sro_n1438;
wire CLOCK_slo__sro_n1439;
wire CLOCK_slo__sro_n1505;
wire CLOCK_slo__sro_n1663;
wire CLOCK_slo__sro_n1507;
wire CLOCK_slo__sro_n1533;
wire CLOCK_slo__sro_n1534;
wire CLOCK_slo__sro_n1535;
wire CLOCK_slo__sro_n1536;
wire CLOCK_slo__sro_n1537;
wire CLOCK_slo__sro_n1604;
wire CLOCK_slo__xsl_n1813;
wire CLOCK_slo__sro_n1592;
wire CLOCK_slo__sro_n1593;
wire CLOCK_slo__sro_n1594;
wire CLOCK_slo__sro_n1595;


INV_X1 i_36 (.ZN (n_34), .A (p_0[30]));
INV_X1 i_35 (.ZN (n_33), .A (p_1[30]));
INV_X1 i_34 (.ZN (n_32), .A (n_30));
INV_X1 slo__sro_c516 (.ZN (slo__sro_n700), .A (n_10));
XOR2_X1 i_32 (.Z (p_2[31]), .A (p_0[31]), .B (slo__sro_n557));
OAI22_X1 i_31 (.ZN (n_0), .A1 (n_34), .A2 (p_1[30]), .B1 (p_0[30]), .B2 (n_33));
XNOR2_X1 i_0 (.ZN (p_2[30]), .A (n_32), .B (n_0));
FA_X1 i_30 (.CO (n_30), .S (p_2[29]), .A (p_0[29]), .B (p_1[29]), .CI (CLOCK_slo__sro_n1534));
OR2_X1 CLOCK_slo__sro_c1176 (.ZN (CLOCK_slo__sro_n1604), .A1 (p_1[14]), .A2 (p_0[14]));
FA_X1 i_28 (.CO (n_28), .S (p_2[27]), .A (p_0[27]), .B (p_1[27]), .CI (n_27));
FA_X1 i_27 (.CO (n_27), .S (p_2[26]), .A (p_0[26]), .B (p_1[26]), .CI (slo__sro_n375));
XNOR2_X1 slo__sro_c326 (.ZN (p_2[21]), .A (slo__sro_n429), .B (CLOCK_slo__xsl_n1812));
INV_X1 slo__sro_c717 (.ZN (slo__sro_n965), .A (n_20));
FA_X1 i_24 (.CO (n_24), .S (p_2[23]), .A (p_0[23]), .B (p_1[23]), .CI (slo__sro_n976));
INV_X1 CLOCK_slo__sro_c988 (.ZN (CLOCK_slo__sro_n1439), .A (n_15));
NOR2_X1 slo__sro_c406 (.ZN (slo__sro_n560), .A1 (n_33), .A2 (p_0[30]));
NAND2_X1 slo__sro_c731 (.ZN (slo__sro_n978), .A1 (slo__sro_n430), .A2 (p_0[22]));
FA_X1 i_20 (.CO (n_20), .S (p_2[19]), .A (p_0[19]), .B (p_1[19]), .CI (slo__sro_n531));
NAND2_X1 slo__sro_c692 (.ZN (slo__sro_n934), .A1 (p_1[24]), .A2 (p_0[24]));
NAND2_X1 slo__sro_c125 (.ZN (slo__sro_n198), .A1 (p_1[16]), .A2 (p_0[16]));
NAND2_X2 slo__sro_c694 (.ZN (n_25), .A1 (slo__sro_n933), .A2 (slo__sro_n934));
NAND2_X1 CLOCK_slo__sro_c1058 (.ZN (CLOCK_slo__sro_n1507), .A1 (p_1[14]), .A2 (p_0[14]));
INV_X1 CLOCK_slo__sro_c1088 (.ZN (CLOCK_slo__sro_n1537), .A (n_28));
INV_X1 slo__sro_c295 (.ZN (slo__sro_n378), .A (p_1[25]));
NOR2_X1 slo__sro_c719 (.ZN (slo__sro_n963), .A1 (opt_ipoPP_5), .A2 (p_0[20]));
FA_X1 i_12 (.CO (n_12), .S (p_2[11]), .A (p_0[11]), .B (p_1[11]), .CI (n_11));
XNOR2_X1 slo__sro_c695 (.ZN (slo__sro_n932), .A (p_1[24]), .B (p_0[24]));
FA_X1 i_10 (.CO (n_10), .S (p_2[9]), .A (p_0[9]), .B (p_1[9]), .CI (n_9));
FA_X1 i_8 (.CO (n_8), .S (p_2[7]), .A (p_0[7]), .B (p_1[7]), .CI (n_7));
FA_X1 i_7 (.CO (n_7), .S (p_2[6]), .A (p_0[6]), .B (p_1[6]), .CI (n_6));
INV_X1 slo__sro_c124 (.ZN (slo__sro_n199), .A (n_16));
FA_X1 i_5 (.CO (n_5), .S (p_2[4]), .A (p_0[4]), .B (p_1[4]), .CI (n_4));
FA_X1 i_4 (.CO (n_4), .S (p_2[3]), .A (p_0[3]), .B (p_1[3]), .CI (n_3));
FA_X1 i_3 (.CO (n_3), .S (p_2[2]), .A (p_0[2]), .B (p_1[2]), .CI (n_2));
FA_X1 i_2 (.CO (n_2), .S (p_2[1]), .A (p_0[1]), .B (p_1[1]), .CI (n_1));
HA_X1 i_1 (.CO (n_1), .S (p_2[0]), .A (p_0[0]), .B (p_1[0]));
INV_X1 slo__sro_c108 (.ZN (slo__sro_n183), .A (n_5));
NAND2_X1 slo__sro_c109 (.ZN (slo__sro_n182), .A1 (p_1[5]), .A2 (p_0[5]));
NOR2_X1 slo__sro_c110 (.ZN (slo__sro_n181), .A1 (p_1[5]), .A2 (p_0[5]));
OAI21_X1 slo__sro_c111 (.ZN (n_6), .A (slo__sro_n182), .B1 (slo__sro_n183), .B2 (slo__sro_n181));
XNOR2_X1 slo__sro_c112 (.ZN (slo__sro_n180), .A (p_1[5]), .B (p_0[5]));
XNOR2_X1 slo__sro_c113 (.ZN (p_2[5]), .A (slo__sro_n180), .B (n_5));
INV_X2 slo__sro_c16 (.ZN (slo__sro_n84), .A (CLOCK_slo__sro_n1663));
NAND2_X1 slo__sro_c17 (.ZN (slo__sro_n83), .A1 (p_1[17]), .A2 (p_0[17]));
NOR2_X2 slo__sro_c18 (.ZN (slo__sro_n82), .A1 (p_1[17]), .A2 (p_0[17]));
OAI21_X2 slo__sro_c19 (.ZN (slo__sro_n81), .A (slo__sro_n83), .B1 (slo__sro_n82), .B2 (slo__sro_n84));
XNOR2_X1 slo__sro_c20 (.ZN (slo__sro_n80), .A (p_1[17]), .B (p_0[17]));
XNOR2_X1 slo__sro_c21 (.ZN (p_2[17]), .A (CLOCK_slo__sro_n1663), .B (slo__sro_n80));
NOR2_X2 slo__sro_c126 (.ZN (slo__sro_n197), .A1 (p_1[16]), .A2 (p_0[16]));
INV_X1 CLOCK_slo__xsl_c1394 (.ZN (CLOCK_slo__xsl_n1813), .A (n_21));
XNOR2_X1 slo__sro_c128 (.ZN (slo__sro_n195), .A (p_1[16]), .B (p_0[16]));
XNOR2_X1 slo__sro_c129 (.ZN (p_2[16]), .A (slo__sro_n195), .B (n_16));
OAI21_X1 slo__sro_c693 (.ZN (slo__sro_n933), .A (n_24), .B1 (p_1[24]), .B2 (p_0[24]));
INV_X1 slo__sro_c405 (.ZN (slo__sro_n561), .A (n_30));
INV_X1 slo__sro_c321 (.ZN (slo__sro_n433), .A (n_21));
NAND2_X1 slo__sro_c322 (.ZN (slo__sro_n432), .A1 (p_0[21]), .A2 (p_1[21]));
NOR2_X1 slo__sro_c323 (.ZN (slo__sro_n431), .A1 (p_1[21]), .A2 (p_0[21]));
OAI21_X2 slo__sro_c324 (.ZN (slo__sro_n430), .A (slo__sro_n432), .B1 (slo__sro_n433), .B2 (slo__sro_n431));
XNOR2_X1 slo__sro_c325 (.ZN (slo__sro_n429), .A (p_1[21]), .B (p_0[21]));
INV_X1 slo__sro_c255 (.ZN (slo__sro_n336), .A (n_13));
NAND2_X1 slo__sro_c256 (.ZN (slo__sro_n335), .A1 (p_0[13]), .A2 (p_1[13]));
NOR2_X1 slo__sro_c257 (.ZN (slo__sro_n334), .A1 (p_1[13]), .A2 (p_0[13]));
OAI21_X1 slo__sro_c258 (.ZN (n_14), .A (slo__sro_n335), .B1 (slo__sro_n336), .B2 (slo__sro_n334));
XNOR2_X1 slo__sro_c259 (.ZN (slo__sro_n333), .A (p_1[13]), .B (p_0[13]));
XNOR2_X1 slo__sro_c260 (.ZN (p_2[13]), .A (n_13), .B (slo__sro_n333));
NAND2_X1 slo__sro_c296 (.ZN (slo__sro_n377), .A1 (n_25), .A2 (p_0[25]));
NOR2_X1 slo__sro_c297 (.ZN (slo__sro_n376), .A1 (n_25), .A2 (p_0[25]));
OAI21_X1 slo__sro_c298 (.ZN (slo__sro_n375), .A (slo__sro_n377), .B1 (slo__sro_n378), .B2 (slo__sro_n376));
XNOR2_X1 slo__sro_c299 (.ZN (slo__sro_n374), .A (n_25), .B (p_0[25]));
XNOR2_X1 slo__sro_c300 (.ZN (p_2[25]), .A (slo__sro_n374), .B (p_1[25]));
NAND2_X1 slo__sro_c407 (.ZN (slo__sro_n559), .A1 (slo__sro_n561), .A2 (slo__sro_n560));
OR2_X1 slo__sro_c408 (.ZN (slo__sro_n558), .A1 (p_1[30]), .A2 (n_34));
OAI21_X1 slo__sro_c409 (.ZN (slo__sro_n557), .A (slo__sro_n559), .B1 (n_32), .B2 (slo__sro_n558));
NAND2_X1 slo__sro_c517 (.ZN (slo__sro_n699), .A1 (p_1[10]), .A2 (p_0[10]));
NOR2_X1 slo__sro_c518 (.ZN (slo__sro_n698), .A1 (p_1[10]), .A2 (p_0[10]));
NAND2_X2 slo__sro_c389 (.ZN (slo__sro_n534), .A1 (p_1[18]), .A2 (p_0[18]));
NAND2_X1 slo__sro_c390 (.ZN (slo__sro_n533), .A1 (slo__sro_n81), .A2 (p_0[18]));
NAND2_X1 slo__sro_c391 (.ZN (slo__sro_n532), .A1 (slo__sro_n81), .A2 (p_1[18]));
NAND3_X1 slo__sro_c392 (.ZN (slo__sro_n531), .A1 (slo__sro_n532), .A2 (slo__sro_n533), .A3 (slo__sro_n534));
XNOR2_X1 slo__sro_c393 (.ZN (slo__sro_n530), .A (slo__sro_n81), .B (p_0[18]));
XNOR2_X2 slo__sro_c394 (.ZN (p_2[18]), .A (slo__sro_n530), .B (p_1[18]));
OAI21_X2 slo__sro_c519 (.ZN (n_11), .A (slo__sro_n699), .B1 (slo__sro_n700), .B2 (slo__sro_n698));
XNOR2_X1 slo__sro_c520 (.ZN (slo__sro_n697), .A (p_1[10]), .B (p_0[10]));
XNOR2_X1 slo__sro_c521 (.ZN (p_2[10]), .A (slo__sro_n697), .B (n_10));
XNOR2_X1 slo__sro_c696 (.ZN (p_2[24]), .A (slo__sro_n932), .B (n_24));
NAND2_X1 slo__sro_c718 (.ZN (slo__sro_n964), .A1 (opt_ipoPP_5), .A2 (p_0[20]));
INV_X1 slo__sro_c676 (.ZN (slo__sro_n918), .A (n_12));
NAND2_X1 slo__sro_c677 (.ZN (slo__sro_n917), .A1 (p_1[12]), .A2 (p_0[12]));
NOR2_X1 slo__sro_c678 (.ZN (slo__sro_n916), .A1 (p_1[12]), .A2 (p_0[12]));
OAI21_X1 slo__sro_c679 (.ZN (n_13), .A (slo__sro_n917), .B1 (slo__sro_n918), .B2 (slo__sro_n916));
XNOR2_X1 slo__sro_c680 (.ZN (slo__sro_n915), .A (p_1[12]), .B (p_0[12]));
XNOR2_X1 slo__sro_c681 (.ZN (p_2[12]), .A (slo__sro_n915), .B (n_12));
OAI21_X2 slo__sro_c720 (.ZN (n_21), .A (slo__sro_n964), .B1 (slo__sro_n965), .B2 (slo__sro_n963));
XNOR2_X1 slo__sro_c721 (.ZN (slo__sro_n962), .A (p_1[20]), .B (p_0[20]));
XNOR2_X1 slo__sro_c722 (.ZN (p_2[20]), .A (slo__sro_n962), .B (n_20));
OAI21_X2 slo__sro_c732 (.ZN (slo__sro_n977), .A (p_1[22]), .B1 (slo__sro_n430), .B2 (p_0[22]));
NAND2_X1 slo__sro_c733 (.ZN (slo__sro_n976), .A1 (slo__sro_n977), .A2 (slo__sro_n978));
XNOR2_X1 slo__sro_c734 (.ZN (slo__sro_n975), .A (slo__sro_n430), .B (p_0[22]));
XNOR2_X1 slo__sro_c735 (.ZN (p_2[22]), .A (slo__sro_n975), .B (p_1[22]));
NAND2_X1 CLOCK_slo__sro_c989 (.ZN (CLOCK_slo__sro_n1438), .A1 (p_1[15]), .A2 (p_0[15]));
NOR2_X1 CLOCK_slo__sro_c990 (.ZN (CLOCK_slo__sro_n1437), .A1 (p_1[15]), .A2 (p_0[15]));
OAI21_X2 CLOCK_slo__sro_c991 (.ZN (n_16), .A (CLOCK_slo__sro_n1438), .B1 (CLOCK_slo__sro_n1439), .B2 (CLOCK_slo__sro_n1437));
XNOR2_X1 CLOCK_slo__sro_c992 (.ZN (CLOCK_slo__sro_n1436), .A (p_1[15]), .B (p_0[15]));
XNOR2_X1 CLOCK_slo__sro_c993 (.ZN (p_2[15]), .A (CLOCK_slo__sro_n1436), .B (n_15));
OAI21_X2 CLOCK_slo__sro_c1240 (.ZN (CLOCK_slo__sro_n1663), .A (slo__sro_n198), .B1 (slo__sro_n199), .B2 (slo__sro_n197));
NAND2_X1 CLOCK_slo__sro_c1060 (.ZN (n_15), .A1 (CLOCK_slo__sro_n1603), .A2 (CLOCK_slo__sro_n1507));
XNOR2_X1 CLOCK_slo__sro_c1061 (.ZN (CLOCK_slo__sro_n1505), .A (p_1[14]), .B (p_0[14]));
XNOR2_X1 CLOCK_slo__sro_c1062 (.ZN (p_2[14]), .A (CLOCK_slo__sro_n1505), .B (n_14));
NAND2_X1 CLOCK_slo__sro_c1089 (.ZN (CLOCK_slo__sro_n1536), .A1 (p_1[28]), .A2 (p_0[28]));
NOR2_X1 CLOCK_slo__sro_c1090 (.ZN (CLOCK_slo__sro_n1535), .A1 (p_1[28]), .A2 (p_0[28]));
OAI21_X1 CLOCK_slo__sro_c1091 (.ZN (CLOCK_slo__sro_n1534), .A (CLOCK_slo__sro_n1536)
    , .B1 (CLOCK_slo__sro_n1535), .B2 (CLOCK_slo__sro_n1537));
XNOR2_X1 CLOCK_slo__sro_c1092 (.ZN (CLOCK_slo__sro_n1533), .A (p_1[28]), .B (p_0[28]));
XNOR2_X1 CLOCK_slo__sro_c1093 (.ZN (p_2[28]), .A (CLOCK_slo__sro_n1533), .B (n_28));
NAND2_X1 CLOCK_slo__sro_c1177 (.ZN (CLOCK_slo__sro_n1603), .A1 (CLOCK_slo__sro_n1604), .A2 (n_14));
INV_X1 CLOCK_slo__xsl_c1395 (.ZN (CLOCK_slo__xsl_n1812), .A (CLOCK_slo__xsl_n1813));
INV_X1 CLOCK_slo__sro_c1162 (.ZN (CLOCK_slo__sro_n1595), .A (n_8));
NAND2_X1 CLOCK_slo__sro_c1163 (.ZN (CLOCK_slo__sro_n1594), .A1 (p_1[8]), .A2 (p_0[8]));
NOR2_X1 CLOCK_slo__sro_c1164 (.ZN (CLOCK_slo__sro_n1593), .A1 (p_1[8]), .A2 (p_0[8]));
OAI21_X1 CLOCK_slo__sro_c1165 (.ZN (n_9), .A (CLOCK_slo__sro_n1594), .B1 (CLOCK_slo__sro_n1595), .B2 (CLOCK_slo__sro_n1593));
XNOR2_X1 CLOCK_slo__sro_c1166 (.ZN (CLOCK_slo__sro_n1592), .A (p_1[8]), .B (p_0[8]));
XNOR2_X1 CLOCK_slo__sro_c1167 (.ZN (p_2[8]), .A (CLOCK_slo__sro_n1592), .B (n_8));

endmodule //datapath__0_222

module datapath__0_221 (Multiplier, p_0, p_1);

output [31:0] p_1;
input [31:0] Multiplier;
input [31:0] p_0;
wire slo__sro_n573;
wire CLOCK_slo__xsl_n1446;
wire slo__sro_n820;
wire n_1;
wire n_2;
wire n_3;
wire n_4;
wire n_5;
wire n_6;
wire n_7;
wire n_8;
wire n_10;
wire n_11;
wire n_12;
wire n_13;
wire slo__sro_n273;
wire n_15;
wire n_18;
wire slo__sro_n779;
wire n_21;
wire n_22;
wire n_23;
wire n_24;
wire n_25;
wire n_28;
wire n_29;
wire n_30;
wire n_32;
wire n_0;
wire n_34;
wire n_33;
wire slo__sro_n59;
wire slo__sro_n60;
wire slo__sro_n61;
wire slo__sro_n62;
wire slo__sro_n72;
wire slo__sro_n73;
wire slo__sro_n74;
wire slo__sro_n75;
wire slo__sro_n91;
wire slo__sro_n92;
wire slo__sro_n93;
wire slo__sro_n94;
wire slo__sro_n106;
wire slo__sro_n107;
wire slo__sro_n108;
wire slo__sro_n109;
wire slo__sro_n119;
wire slo__sro_n120;
wire slo__sro_n121;
wire slo__sro_n122;
wire slo__sro_n136;
wire slo__sro_n137;
wire slo__sro_n138;
wire slo__sro_n139;
wire slo__sro_n153;
wire slo__sro_n154;
wire slo__sro_n155;
wire slo__sro_n156;
wire slo__sro_n168;
wire slo__sro_n169;
wire slo__sro_n170;
wire CLOCK_slo__sro_n1313;
wire slo__sro_n179;
wire slo__sro_n180;
wire slo__sro_n181;
wire slo__sro_n182;
wire slo__sro_n183;
wire slo__sro_n216;
wire slo__sro_n217;
wire slo__sro_n218;
wire slo__sro_n231;
wire slo__sro_n233;
wire slo__sro_n274;
wire slo__sro_n275;
wire slo__sro_n276;
wire slo__sro_n277;
wire slo__sro_n291;
wire slo__sro_n292;
wire slo__sro_n293;
wire slo__sro_n294;
wire slo__sro_n375;
wire CLOCK_slo__mro_n1432;
wire slo__sro_n331;
wire slo__sro_n332;
wire slo__sro_n376;
wire slo__sro_n377;
wire slo__sro_n378;
wire slo__sro_n379;
wire slo__sro_n459;
wire slo__sro_n460;
wire slo__sro_n461;
wire slo__sro_n574;
wire slo__sro_n575;
wire slo__sro_n576;
wire slo__sro_n577;
wire slo__sro_n780;
wire slo__sro_n781;
wire slo__sro_n782;
wire slo__mro_n807;
wire slo__sro_n821;
wire slo__sro_n822;
wire slo__sro_n823;
wire slo__sro_n824;
wire slo__sro_n861;
wire slo__sro_n862;
wire slo__sro_n863;
wire slo__sro_n1132;
wire slo__sro_n1133;
wire slo__sro_n1134;
wire slo__sro_n1135;
wire slo__sro_n1136;
wire CLOCK_slo__mro_n1283;
wire CLOCK_slo__sro_n1314;
wire CLOCK_slo__sro_n1315;
wire CLOCK_slo__sro_n1316;
wire CLOCK_slo__sro_n1345;
wire CLOCK_slo__sro_n1346;
wire CLOCK_slo__sro_n1347;
wire CLOCK_slo__sro_n1348;
wire CLOCK_slo__sro_n1357;
wire CLOCK_slo__sro_n1358;
wire CLOCK_slo__sro_n1359;
wire CLOCK_slo__sro_n1360;
wire CLOCK_slo__mro_n1421;
wire CLOCK_slo__sro_n1517;
wire CLOCK_slo__sro_n1518;
wire CLOCK_slo__sro_n1519;


INV_X1 i_36 (.ZN (n_34), .A (Multiplier[30]));
INV_X2 i_35 (.ZN (n_33), .A (p_0[30]));
INV_X1 i_34 (.ZN (n_32), .A (n_30));
INV_X2 slo__sro_c401 (.ZN (slo__sro_n577), .A (n_18));
XOR2_X1 i_32 (.Z (p_1[31]), .A (Multiplier[31]), .B (slo__sro_n273));
OAI22_X1 i_31 (.ZN (n_0), .A1 (n_34), .A2 (p_0[30]), .B1 (n_33), .B2 (Multiplier[30]));
XNOR2_X1 i_0 (.ZN (p_1[30]), .A (n_32), .B (n_0));
FA_X1 i_30 (.CO (n_30), .S (p_1[29]), .A (Multiplier[29]), .B (p_0[29]), .CI (n_29));
XNOR2_X2 slo__mro_c539 (.ZN (slo__mro_n807), .A (p_0[13]), .B (Multiplier[13]));
INV_X1 CLOCK_slo__sro_c913 (.ZN (CLOCK_slo__sro_n1348), .A (p_0[13]));
NAND2_X1 slo__sro_c402 (.ZN (slo__sro_n576), .A1 (p_0[18]), .A2 (Multiplier[18]));
INV_X1 slo__sro_c151 (.ZN (slo__sro_n218), .A (n_3));
NOR2_X2 slo__sro_c263 (.ZN (slo__sro_n377), .A1 (p_0[19]), .A2 (Multiplier[19]));
XNOR2_X2 CLOCK_slo__mro_c998 (.ZN (CLOCK_slo__mro_n1421), .A (p_0[24]), .B (Multiplier[24]));
INV_X1 slo__sro_c57 (.ZN (slo__sro_n122), .A (n_10));
INV_X2 slo__sro_c261 (.ZN (slo__sro_n379), .A (slo__sro_n574));
FA_X1 i_21 (.CO (n_21), .S (p_1[20]), .A (Multiplier[20]), .B (p_0[20]), .CI (slo__sro_n376));
XNOR2_X1 slo__sro_c298 (.ZN (p_1[25]), .A (p_0[25]), .B (slo__sro_n179));
NAND2_X1 slo__sro_c520 (.ZN (slo__sro_n781), .A1 (p_0[28]), .A2 (Multiplier[28]));
NAND2_X1 slo__sro_c582 (.ZN (slo__sro_n863), .A1 (p_0[9]), .A2 (Multiplier[9]));
NAND2_X1 slo__sro_c31 (.ZN (slo__sro_n94), .A1 (p_0[15]), .A2 (Multiplier[15]));
INV_X1 slo__sro_c43 (.ZN (slo__sro_n109), .A (n_22));
NAND2_X1 CLOCK_slo__sro_c1193 (.ZN (slo__sro_n108), .A1 (p_0[22]), .A2 (Multiplier[22]));
INV_X1 slo__sro_c185 (.ZN (slo__sro_n277), .A (n_30));
FA_X1 i_13 (.CO (n_13), .S (p_1[12]), .A (Multiplier[12]), .B (p_0[12]), .CI (n_12));
INV_X2 slo__sro_c115 (.ZN (slo__sro_n183), .A (p_0[25]));
INV_X1 slo__sro_c73 (.ZN (slo__sro_n139), .A (n_5));
NAND2_X1 slo__sro_c728 (.ZN (slo__sro_n1135), .A1 (p_0[8]), .A2 (Multiplier[8]));
XNOR2_X2 CLOCK_slo__mro_c844 (.ZN (CLOCK_slo__mro_n1283), .A (slo__sro_n180), .B (Multiplier[26]));
FA_X1 i_8 (.CO (n_8), .S (p_1[7]), .A (Multiplier[7]), .B (p_0[7]), .CI (n_7));
NAND2_X1 CLOCK_slo__sro_c1104 (.ZN (CLOCK_slo__sro_n1519), .A1 (p_0[14]), .A2 (Multiplier[14]));
INV_X1 slo__sro_c89 (.ZN (slo__sro_n156), .A (n_4));
NAND2_X1 slo__sro_c103 (.ZN (slo__sro_n170), .A1 (n_11), .A2 (Multiplier[11]));
NAND2_X1 slo__sro_c165 (.ZN (slo__sro_n233), .A1 (Multiplier[13]), .A2 (p_0[13]));
FA_X1 i_3 (.CO (n_3), .S (p_1[2]), .A (Multiplier[2]), .B (p_0[2]), .CI (n_2));
FA_X1 i_2 (.CO (n_2), .S (p_1[1]), .A (Multiplier[1]), .B (p_0[1]), .CI (n_1));
HA_X1 i_1 (.CO (n_1), .S (p_1[0]), .A (Multiplier[0]), .B (p_0[0]));
INV_X1 slo__sro_c1 (.ZN (slo__sro_n62), .A (n_6));
NAND2_X1 slo__sro_c2 (.ZN (slo__sro_n61), .A1 (p_0[6]), .A2 (Multiplier[6]));
NOR2_X1 slo__sro_c3 (.ZN (slo__sro_n60), .A1 (p_0[6]), .A2 (Multiplier[6]));
OAI21_X1 slo__sro_c4 (.ZN (n_7), .A (slo__sro_n61), .B1 (slo__sro_n60), .B2 (slo__sro_n62));
XNOR2_X1 slo__sro_c5 (.ZN (slo__sro_n59), .A (p_0[6]), .B (Multiplier[6]));
XNOR2_X1 slo__sro_c6 (.ZN (p_1[6]), .A (slo__sro_n59), .B (n_6));
NAND2_X1 slo__sro_c16 (.ZN (slo__sro_n75), .A1 (p_0[16]), .A2 (Multiplier[16]));
NOR2_X2 slo__sro_c17 (.ZN (slo__sro_n74), .A1 (p_0[16]), .A2 (Multiplier[16]));
OAI21_X1 slo__sro_c18 (.ZN (slo__sro_n73), .A (slo__sro_n75), .B1 (slo__sro_n74), .B2 (slo__sro_n92));
XNOR2_X1 slo__sro_c19 (.ZN (slo__sro_n72), .A (p_0[16]), .B (Multiplier[16]));
XNOR2_X1 slo__sro_c20 (.ZN (p_1[16]), .A (slo__sro_n72), .B (CLOCK_slo__xsl_n1446));
OAI21_X1 slo__sro_c32 (.ZN (slo__sro_n93), .A (n_15), .B1 (p_0[15]), .B2 (Multiplier[15]));
NAND2_X1 CLOCK_slo__sro_c1106 (.ZN (n_15), .A1 (CLOCK_slo__sro_n1518), .A2 (CLOCK_slo__sro_n1519));
XNOR2_X1 slo__sro_c34 (.ZN (slo__sro_n91), .A (p_0[15]), .B (Multiplier[15]));
XNOR2_X1 slo__sro_c35 (.ZN (p_1[15]), .A (slo__sro_n91), .B (n_15));
NOR2_X2 slo__sro_c45 (.ZN (slo__sro_n107), .A1 (p_0[22]), .A2 (Multiplier[22]));
INV_X1 slo__sro_c727 (.ZN (slo__sro_n1136), .A (n_8));
XNOR2_X2 slo__sro_c47 (.ZN (slo__sro_n106), .A (p_0[22]), .B (Multiplier[22]));
XNOR2_X2 slo__sro_c48 (.ZN (p_1[22]), .A (slo__sro_n106), .B (n_22));
NAND2_X1 slo__sro_c58 (.ZN (slo__sro_n121), .A1 (p_0[10]), .A2 (Multiplier[10]));
NOR2_X2 slo__sro_c59 (.ZN (slo__sro_n120), .A1 (p_0[10]), .A2 (Multiplier[10]));
OAI21_X2 slo__sro_c60 (.ZN (n_11), .A (slo__sro_n121), .B1 (slo__sro_n120), .B2 (slo__sro_n122));
XNOR2_X2 slo__sro_c61 (.ZN (slo__sro_n119), .A (p_0[10]), .B (Multiplier[10]));
XNOR2_X1 slo__sro_c62 (.ZN (p_1[10]), .A (slo__sro_n119), .B (n_10));
NAND2_X1 slo__sro_c74 (.ZN (slo__sro_n138), .A1 (p_0[5]), .A2 (Multiplier[5]));
NOR2_X1 slo__sro_c75 (.ZN (slo__sro_n137), .A1 (p_0[5]), .A2 (Multiplier[5]));
OAI21_X1 slo__sro_c76 (.ZN (n_6), .A (slo__sro_n138), .B1 (slo__sro_n139), .B2 (slo__sro_n137));
XNOR2_X2 slo__sro_c77 (.ZN (slo__sro_n136), .A (p_0[5]), .B (Multiplier[5]));
XNOR2_X1 slo__sro_c78 (.ZN (p_1[5]), .A (slo__sro_n136), .B (n_5));
NAND2_X1 slo__sro_c90 (.ZN (slo__sro_n155), .A1 (p_0[4]), .A2 (Multiplier[4]));
NOR2_X1 slo__sro_c91 (.ZN (slo__sro_n154), .A1 (p_0[4]), .A2 (Multiplier[4]));
OAI21_X1 slo__sro_c92 (.ZN (n_5), .A (slo__sro_n155), .B1 (slo__sro_n154), .B2 (slo__sro_n156));
XNOR2_X1 slo__sro_c93 (.ZN (slo__sro_n153), .A (p_0[4]), .B (Multiplier[4]));
XNOR2_X1 slo__sro_c94 (.ZN (p_1[4]), .A (slo__sro_n153), .B (n_4));
OAI21_X2 slo__sro_c104 (.ZN (slo__sro_n169), .A (p_0[11]), .B1 (n_11), .B2 (Multiplier[11]));
NAND2_X1 slo__sro_c105 (.ZN (n_12), .A1 (slo__sro_n169), .A2 (slo__sro_n170));
XNOR2_X1 slo__sro_c106 (.ZN (slo__sro_n168), .A (n_11), .B (Multiplier[11]));
XNOR2_X1 slo__sro_c107 (.ZN (p_1[11]), .A (slo__sro_n168), .B (p_0[11]));
NAND2_X1 slo__sro_c116 (.ZN (slo__sro_n182), .A1 (n_25), .A2 (Multiplier[25]));
NOR2_X1 slo__sro_c117 (.ZN (slo__sro_n181), .A1 (n_25), .A2 (Multiplier[25]));
OAI21_X2 slo__sro_c118 (.ZN (slo__sro_n180), .A (slo__sro_n182), .B1 (slo__sro_n183), .B2 (slo__sro_n181));
XNOR2_X1 slo__sro_c119 (.ZN (slo__sro_n179), .A (n_25), .B (Multiplier[25]));
NAND2_X1 slo__sro_c323 (.ZN (slo__sro_n461), .A1 (p_0[26]), .A2 (Multiplier[26]));
NAND2_X1 slo__sro_c152 (.ZN (slo__sro_n217), .A1 (p_0[3]), .A2 (Multiplier[3]));
NOR2_X1 slo__sro_c153 (.ZN (slo__sro_n216), .A1 (p_0[3]), .A2 (Multiplier[3]));
OAI21_X1 slo__sro_c154 (.ZN (n_4), .A (slo__sro_n217), .B1 (slo__sro_n216), .B2 (slo__sro_n218));
BUF_X4 CLOCK_slo__sro_c923 (.Z (CLOCK_slo__sro_n1360), .A (n_23));
NAND2_X1 slo__sro_c167 (.ZN (slo__sro_n231), .A1 (CLOCK_slo__sro_n1345), .A2 (slo__sro_n233));
BUF_X4 slo__sro_c549 (.Z (slo__sro_n824), .A (slo__sro_n73));
NAND2_X1 slo__sro_c550 (.ZN (slo__sro_n823), .A1 (p_0[17]), .A2 (Multiplier[17]));
NOR2_X1 slo__sro_c186 (.ZN (slo__sro_n276), .A1 (n_33), .A2 (Multiplier[30]));
NAND2_X1 slo__sro_c187 (.ZN (slo__sro_n275), .A1 (slo__sro_n276), .A2 (slo__sro_n277));
OR2_X1 slo__sro_c188 (.ZN (slo__sro_n274), .A1 (p_0[30]), .A2 (n_34));
OAI21_X1 slo__sro_c189 (.ZN (slo__sro_n273), .A (slo__sro_n275), .B1 (n_32), .B2 (slo__sro_n274));
INV_X1 slo__sro_c201 (.ZN (slo__sro_n294), .A (n_21));
NAND2_X1 slo__sro_c202 (.ZN (slo__sro_n293), .A1 (p_0[21]), .A2 (Multiplier[21]));
NOR2_X1 slo__sro_c203 (.ZN (slo__sro_n292), .A1 (p_0[21]), .A2 (Multiplier[21]));
OAI21_X2 slo__sro_c204 (.ZN (n_22), .A (slo__sro_n293), .B1 (slo__sro_n294), .B2 (slo__sro_n292));
XNOR2_X1 slo__sro_c205 (.ZN (slo__sro_n291), .A (p_0[21]), .B (Multiplier[21]));
XNOR2_X1 slo__sro_c206 (.ZN (p_1[21]), .A (slo__sro_n291), .B (n_21));
NAND2_X1 slo__sro_c262 (.ZN (slo__sro_n378), .A1 (p_0[19]), .A2 (Multiplier[19]));
NAND2_X1 slo__sro_c231 (.ZN (slo__sro_n332), .A1 (p_0[24]), .A2 (Multiplier[24]));
OAI21_X2 slo__sro_c232 (.ZN (slo__sro_n331), .A (n_24), .B1 (p_0[24]), .B2 (Multiplier[24]));
NAND2_X2 slo__sro_c233 (.ZN (n_25), .A1 (slo__sro_n331), .A2 (slo__sro_n332));
XNOR2_X2 CLOCK_slo__mro_c1006 (.ZN (CLOCK_slo__mro_n1432), .A (p_0[3]), .B (Multiplier[3]));
XNOR2_X1 CLOCK_slo__mro_c1007 (.ZN (p_1[3]), .A (CLOCK_slo__mro_n1432), .B (n_3));
OAI21_X2 slo__sro_c264 (.ZN (slo__sro_n376), .A (slo__sro_n378), .B1 (slo__sro_n379), .B2 (slo__sro_n377));
XNOR2_X1 slo__sro_c265 (.ZN (slo__sro_n375), .A (p_0[19]), .B (Multiplier[19]));
XNOR2_X1 slo__sro_c266 (.ZN (p_1[19]), .A (slo__sro_n375), .B (slo__sro_n574));
OAI21_X1 slo__sro_c324 (.ZN (slo__sro_n460), .A (slo__sro_n180), .B1 (p_0[26]), .B2 (Multiplier[26]));
NAND2_X2 slo__sro_c325 (.ZN (slo__sro_n459), .A1 (slo__sro_n460), .A2 (slo__sro_n461));
NAND2_X2 CLOCK_slo__sro_c879 (.ZN (CLOCK_slo__sro_n1316), .A1 (p_0[27]), .A2 (Multiplier[27]));
NAND2_X1 CLOCK_slo__sro_c880 (.ZN (CLOCK_slo__sro_n1315), .A1 (slo__sro_n459), .A2 (Multiplier[27]));
NOR2_X2 slo__sro_c403 (.ZN (slo__sro_n575), .A1 (p_0[18]), .A2 (Multiplier[18]));
INV_X1 slo__sro_c519 (.ZN (slo__sro_n782), .A (n_28));
OAI21_X1 CLOCK_slo__sro_c1105 (.ZN (CLOCK_slo__sro_n1518), .A (slo__sro_n231), .B1 (p_0[14]), .B2 (Multiplier[14]));
XNOR2_X1 slo__sro_c405 (.ZN (slo__sro_n573), .A (p_0[18]), .B (Multiplier[18]));
XNOR2_X1 slo__sro_c406 (.ZN (p_1[18]), .A (n_18), .B (slo__sro_n573));
NOR2_X2 slo__sro_c521 (.ZN (slo__sro_n780), .A1 (p_0[28]), .A2 (Multiplier[28]));
OAI21_X2 slo__sro_c522 (.ZN (n_29), .A (slo__sro_n781), .B1 (slo__sro_n780), .B2 (slo__sro_n782));
XNOR2_X1 slo__sro_c523 (.ZN (slo__sro_n779), .A (p_0[28]), .B (Multiplier[28]));
XNOR2_X1 slo__sro_c524 (.ZN (p_1[28]), .A (slo__sro_n779), .B (n_28));
XNOR2_X2 slo__mro_c540 (.ZN (p_1[13]), .A (n_13), .B (slo__mro_n807));
NAND2_X2 slo__sro_c551 (.ZN (slo__sro_n822), .A1 (slo__sro_n824), .A2 (Multiplier[17]));
NAND2_X2 slo__sro_c552 (.ZN (slo__sro_n821), .A1 (slo__sro_n824), .A2 (p_0[17]));
NAND3_X4 slo__sro_c553 (.ZN (n_18), .A1 (slo__sro_n822), .A2 (slo__sro_n821), .A3 (slo__sro_n823));
XNOR2_X2 slo__sro_c554 (.ZN (slo__sro_n820), .A (p_0[17]), .B (Multiplier[17]));
XNOR2_X2 slo__sro_c555 (.ZN (p_1[17]), .A (slo__sro_n820), .B (slo__sro_n824));
OAI21_X1 slo__sro_c583 (.ZN (slo__sro_n862), .A (slo__sro_n1133), .B1 (p_0[9]), .B2 (Multiplier[9]));
NAND2_X1 slo__sro_c584 (.ZN (n_10), .A1 (slo__sro_n862), .A2 (slo__sro_n863));
XNOR2_X1 slo__sro_c585 (.ZN (slo__sro_n861), .A (p_0[9]), .B (Multiplier[9]));
XNOR2_X1 slo__sro_c586 (.ZN (p_1[9]), .A (slo__sro_n861), .B (slo__sro_n1133));
NOR2_X1 slo__sro_c729 (.ZN (slo__sro_n1134), .A1 (p_0[8]), .A2 (Multiplier[8]));
OAI21_X1 slo__sro_c646 (.ZN (n_23), .A (slo__sro_n108), .B1 (slo__sro_n107), .B2 (slo__sro_n109));
OAI21_X1 slo__sro_c730 (.ZN (slo__sro_n1133), .A (slo__sro_n1135), .B1 (slo__sro_n1136), .B2 (slo__sro_n1134));
XNOR2_X2 slo__sro_c731 (.ZN (slo__sro_n1132), .A (p_0[8]), .B (Multiplier[8]));
XNOR2_X1 slo__sro_c732 (.ZN (p_1[8]), .A (slo__sro_n1132), .B (n_8));
XNOR2_X2 CLOCK_slo__mro_c845 (.ZN (p_1[26]), .A (CLOCK_slo__mro_n1283), .B (p_0[26]));
NAND2_X1 CLOCK_slo__sro_c881 (.ZN (CLOCK_slo__sro_n1314), .A1 (slo__sro_n459), .A2 (p_0[27]));
NAND3_X4 CLOCK_slo__sro_c882 (.ZN (n_28), .A1 (CLOCK_slo__sro_n1315), .A2 (CLOCK_slo__sro_n1314), .A3 (CLOCK_slo__sro_n1316));
XNOR2_X1 CLOCK_slo__sro_c883 (.ZN (CLOCK_slo__sro_n1313), .A (p_0[27]), .B (Multiplier[27]));
XNOR2_X1 CLOCK_slo__sro_c884 (.ZN (p_1[27]), .A (CLOCK_slo__sro_n1313), .B (slo__sro_n459));
INV_X1 CLOCK_slo__sro_c914 (.ZN (CLOCK_slo__sro_n1347), .A (Multiplier[13]));
NAND2_X1 CLOCK_slo__sro_c915 (.ZN (CLOCK_slo__sro_n1346), .A1 (CLOCK_slo__sro_n1348), .A2 (CLOCK_slo__sro_n1347));
NAND2_X1 CLOCK_slo__sro_c916 (.ZN (CLOCK_slo__sro_n1345), .A1 (n_13), .A2 (CLOCK_slo__sro_n1346));
NAND2_X1 CLOCK_slo__sro_c924 (.ZN (CLOCK_slo__sro_n1359), .A1 (CLOCK_slo__sro_n1360), .A2 (Multiplier[23]));
AOI22_X4 CLOCK_slo__sro_c925 (.ZN (CLOCK_slo__sro_n1358), .A1 (CLOCK_slo__sro_n1360)
    , .A2 (p_0[23]), .B1 (p_0[23]), .B2 (Multiplier[23]));
NAND2_X4 CLOCK_slo__sro_c926 (.ZN (n_24), .A1 (CLOCK_slo__sro_n1358), .A2 (CLOCK_slo__sro_n1359));
XNOR2_X2 CLOCK_slo__sro_c927 (.ZN (CLOCK_slo__sro_n1357), .A (p_0[23]), .B (Multiplier[23]));
XNOR2_X2 CLOCK_slo__sro_c928 (.ZN (p_1[23]), .A (CLOCK_slo__sro_n1357), .B (CLOCK_slo__sro_n1360));
XNOR2_X2 CLOCK_slo__mro_c999 (.ZN (p_1[24]), .A (CLOCK_slo__mro_n1421), .B (n_24));
OAI21_X4 CLOCK_slo__sro_c1094 (.ZN (slo__sro_n574), .A (slo__sro_n576), .B1 (slo__sro_n577), .B2 (slo__sro_n575));
INV_X1 CLOCK_slo__xsl_c1023 (.ZN (CLOCK_slo__xsl_n1446), .A (slo__sro_n92));
AND2_X1 CLOCK_slo__xsl_c1026 (.ZN (slo__sro_n92), .A1 (slo__sro_n93), .A2 (slo__sro_n94));
XNOR2_X1 CLOCK_slo__sro_c1107 (.ZN (CLOCK_slo__sro_n1517), .A (p_0[14]), .B (Multiplier[14]));
XNOR2_X1 CLOCK_slo__sro_c1108 (.ZN (p_1[14]), .A (CLOCK_slo__sro_n1517), .B (slo__sro_n231));

endmodule //datapath__0_221

module datapath__0_217 (p_0, p_1, p_2);

output [31:0] p_2;
input [31:0] p_0;
input [31:0] p_1;
wire n_1;
wire n_2;
wire n_4;
wire n_8;
wire n_9;
wire n_10;
wire n_11;
wire n_12;
wire n_14;
wire n_15;
wire CLOCK_slo__sro_n1532;
wire n_17;
wire n_18;
wire slo__sro_n267;
wire n_20;
wire n_21;
wire n_22;
wire n_24;
wire n_25;
wire n_26;
wire n_27;
wire n_28;
wire n_29;
wire n_30;
wire n_32;
wire n_0;
wire n_34;
wire n_33;
wire slo__sro_n63;
wire slo__sro_n64;
wire slo__sro_n65;
wire slo__sro_n66;
wire slo__sro_n472;
wire slo__sro_n100;
wire slo__sro_n101;
wire slo__sro_n102;
wire slo__sro_n103;
wire slo__sro_n104;
wire slo__sro_n216;
wire slo__sro_n217;
wire slo__sro_n218;
wire slo__sro_n170;
wire slo__sro_n171;
wire slo__sro_n172;
wire slo__sro_n173;
wire slo__sro_n174;
wire slo__sro_n202;
wire slo__sro_n203;
wire slo__sro_n204;
wire slo__sro_n205;
wire slo__sro_n268;
wire slo__sro_n269;
wire slo__sro_n270;
wire slo__sro_n271;
wire slo__sro_n319;
wire slo__sro_n320;
wire slo__sro_n321;
wire slo__sro_n322;
wire slo__n339;
wire CLOCK_slo__sro_n2059;
wire slo__sro_n474;
wire slo__sro_n481;
wire slo__sro_n482;
wire slo__sro_n483;
wire slo__sro_n484;
wire slo__sro_n485;
wire slo__sro_n604;
wire slo__sro_n403;
wire slo__sro_n404;
wire slo__sro_n405;
wire CLOCK_slo__sro_n1216;
wire slo__sro_n605;
wire slo__sro_n606;
wire slo__sro_n607;
wire slo__sro_n608;
wire slo__mro_n638;
wire slo__n869;
wire CLOCK_slo__sro_n1217;
wire slo__sro_n996;
wire slo__sro_n997;
wire slo__sro_n998;
wire slo__sro_n999;
wire CLOCK_slo__sro_n1218;
wire CLOCK_slo__sro_n1219;
wire CLOCK_slo__sro_n1220;
wire CLOCK_slo__sro_n1325;
wire CLOCK_slo__sro_n1326;
wire CLOCK_slo__sro_n1327;
wire CLOCK_slo__sro_n1328;
wire CLOCK_slo__sro_n1329;
wire CLOCK_slo__sro_n1533;
wire CLOCK_slo__sro_n1534;
wire CLOCK_slo__sro_n1535;
wire CLOCK_slo__sro_n1385;
wire CLOCK_slo__sro_n1386;
wire CLOCK_slo__sro_n1387;
wire CLOCK_slo__sro_n1388;


INV_X1 i_36 (.ZN (n_34), .A (p_0[30]));
INV_X1 i_35 (.ZN (n_33), .A (p_1[30]));
INV_X1 i_34 (.ZN (n_32), .A (n_30));
INV_X1 slo__sro_c436 (.ZN (slo__sro_n608), .A (slo__sro_n216));
XOR2_X1 i_32 (.Z (p_2[31]), .A (p_0[31]), .B (slo__sro_n481));
OAI22_X1 i_31 (.ZN (n_0), .A1 (n_34), .A2 (p_1[30]), .B1 (p_0[30]), .B2 (n_33));
XNOR2_X1 i_0 (.ZN (p_2[30]), .A (n_32), .B (n_0));
FA_X1 i_30 (.CO (n_30), .S (p_2[29]), .A (p_0[29]), .B (p_1[29]), .CI (n_29));
XNOR2_X2 slo__sro_c321 (.ZN (p_2[6]), .A (slo__sro_n605), .B (slo__sro_n100));
FA_X1 i_28 (.CO (n_28), .S (p_2[27]), .A (p_0[27]), .B (p_1[27]), .CI (n_27));
FA_X1 i_27 (.CO (n_27), .S (p_2[26]), .A (p_0[26]), .B (p_1[26]), .CI (n_26));
FA_X1 i_26 (.CO (n_26), .S (p_2[25]), .A (p_0[25]), .B (p_1[25]), .CI (n_25));
FA_X1 i_24 (.CO (n_24), .S (p_2[23]), .A (p_0[23]), .B (p_1[23]), .CI (CLOCK_slo__sro_n2059));
XNOR2_X1 CLOCK_slo__sro_c832 (.ZN (CLOCK_slo__sro_n1216), .A (p_1[2]), .B (p_0[2]));
INV_X1 slo__sro_c373 (.ZN (slo__sro_n485), .A (n_30));
FA_X1 i_21 (.CO (n_21), .S (p_2[20]), .A (p_0[20]), .B (p_1[20]), .CI (n_20));
XNOR2_X1 slo__sro_c440 (.ZN (slo__sro_n604), .A (p_1[5]), .B (p_0[5]));
INV_X1 slo__sro_c136 (.ZN (slo__sro_n205), .A (n_11));
INV_X1 slo__sro_c41 (.ZN (slo__sro_n104), .A (slo__sro_n605));
FA_X1 i_17 (.CO (n_17), .S (p_2[16]), .A (p_0[16]), .B (p_1[16]), .CI (CLOCK_slo__sro_n1326));
FA_X1 i_15 (.CO (n_15), .S (p_2[14]), .A (p_0[14]), .B (p_1[14]), .CI (n_14));
FA_X1 i_14 (.CO (n_14), .S (p_2[13]), .A (p_0[13]), .B (p_1[13]), .CI (slo__sro_n268));
NAND2_X1 slo__sro_c361 (.ZN (slo__sro_n474), .A1 (p_1[21]), .A2 (p_0[21]));
NOR2_X1 slo__sro_c203 (.ZN (slo__sro_n269), .A1 (p_1[12]), .A2 (p_0[12]));
FA_X1 i_11 (.CO (n_11), .S (p_2[10]), .A (p_0[10]), .B (p_1[10]), .CI (n_10));
FA_X1 i_10 (.CO (n_10), .S (p_2[9]), .A (p_0[9]), .B (p_1[9]), .CI (n_9));
FA_X1 i_9 (.CO (n_9), .S (p_2[8]), .A (p_0[8]), .B (p_1[8]), .CI (n_8));
FA_X1 i_8 (.CO (n_8), .S (p_2[7]), .A (p_0[7]), .B (p_1[7]), .CI (slo__sro_n101));
NAND2_X1 slo__sro_c150 (.ZN (slo__sro_n218), .A1 (n_4), .A2 (p_0[4]));
XNOR2_X1 slo__mro_c461 (.ZN (slo__mro_n638), .A (p_1[4]), .B (p_0[4]));
INV_X2 slo__sro_c201 (.ZN (slo__sro_n271), .A (n_12));
FA_X1 i_4 (.CO (n_4), .S (p_2[3]), .A (p_0[3]), .B (p_1[3]), .CI (CLOCK_slo__sro_n1217));
INV_X2 CLOCK_slo__sro_c933 (.ZN (CLOCK_slo__sro_n1329), .A (n_15));
FA_X1 i_2 (.CO (n_2), .S (p_2[1]), .A (p_0[1]), .B (p_1[1]), .CI (n_1));
HA_X1 i_1 (.CO (n_1), .S (p_2[0]), .A (p_0[0]), .B (p_1[0]));
INV_X1 slo__sro_c1 (.ZN (slo__sro_n66), .A (n_17));
NAND2_X1 slo__sro_c2 (.ZN (slo__sro_n65), .A1 (p_1[17]), .A2 (p_0[17]));
NOR2_X1 slo__sro_c3 (.ZN (slo__sro_n64), .A1 (p_1[17]), .A2 (p_0[17]));
OAI21_X1 slo__sro_c4 (.ZN (n_18), .A (slo__sro_n65), .B1 (slo__sro_n66), .B2 (slo__sro_n64));
XNOR2_X1 slo__sro_c5 (.ZN (slo__sro_n63), .A (p_1[17]), .B (p_0[17]));
XNOR2_X1 slo__sro_c6 (.ZN (p_2[17]), .A (n_17), .B (slo__sro_n63));
NAND2_X1 slo__sro_c42 (.ZN (slo__sro_n103), .A1 (p_1[6]), .A2 (p_0[6]));
NOR2_X1 slo__sro_c43 (.ZN (slo__sro_n102), .A1 (p_1[6]), .A2 (p_0[6]));
OAI21_X1 slo__sro_c44 (.ZN (slo__sro_n101), .A (slo__sro_n103), .B1 (slo__sro_n102), .B2 (slo__sro_n104));
XNOR2_X2 slo__sro_c45 (.ZN (slo__sro_n100), .A (p_1[6]), .B (p_0[6]));
OAI21_X1 CLOCK_slo__sro_c1690 (.ZN (CLOCK_slo__sro_n2059), .A (slo__sro_n998), .B1 (slo__sro_n999), .B2 (slo__sro_n997));
OAI21_X1 slo__sro_c151 (.ZN (slo__sro_n217), .A (p_1[4]), .B1 (n_4), .B2 (p_0[4]));
NAND2_X1 slo__sro_c152 (.ZN (slo__sro_n216), .A1 (slo__sro_n218), .A2 (slo__sro_n217));
NAND2_X1 slo__sro_c202 (.ZN (slo__sro_n270), .A1 (p_1[12]), .A2 (p_0[12]));
INV_X1 slo__sro_c109 (.ZN (slo__sro_n174), .A (slo__n339));
NAND2_X1 slo__sro_c110 (.ZN (slo__sro_n173), .A1 (p_1[18]), .A2 (p_0[18]));
NOR2_X1 slo__sro_c111 (.ZN (slo__sro_n172), .A1 (p_1[18]), .A2 (p_0[18]));
OAI21_X2 slo__sro_c112 (.ZN (slo__sro_n171), .A (slo__sro_n173), .B1 (slo__sro_n174), .B2 (slo__sro_n172));
XNOR2_X1 slo__sro_c113 (.ZN (slo__sro_n170), .A (p_1[18]), .B (p_0[18]));
XNOR2_X1 slo__sro_c114 (.ZN (p_2[18]), .A (n_18), .B (slo__sro_n170));
NAND2_X1 slo__sro_c137 (.ZN (slo__sro_n204), .A1 (p_1[11]), .A2 (p_0[11]));
NOR2_X1 slo__sro_c138 (.ZN (slo__sro_n203), .A1 (p_1[11]), .A2 (p_0[11]));
INV_X1 CLOCK_slo__sro_c1129 (.ZN (CLOCK_slo__sro_n1535), .A (p_1[21]));
XNOR2_X1 slo__sro_c140 (.ZN (slo__sro_n202), .A (p_1[11]), .B (p_0[11]));
XNOR2_X1 slo__sro_c141 (.ZN (p_2[11]), .A (slo__sro_n202), .B (n_11));
OAI21_X1 slo__sro_c204 (.ZN (slo__sro_n268), .A (slo__sro_n270), .B1 (slo__sro_n271), .B2 (slo__sro_n269));
XNOR2_X1 slo__sro_c205 (.ZN (slo__sro_n267), .A (p_1[12]), .B (p_0[12]));
XNOR2_X1 slo__sro_c206 (.ZN (p_2[12]), .A (slo__sro_n267), .B (n_12));
INV_X1 slo__sro_c227 (.ZN (slo__sro_n322), .A (n_28));
NAND2_X1 slo__sro_c228 (.ZN (slo__sro_n321), .A1 (p_1[28]), .A2 (p_0[28]));
NOR2_X1 slo__sro_c229 (.ZN (slo__sro_n320), .A1 (p_1[28]), .A2 (p_0[28]));
OAI21_X1 slo__sro_c230 (.ZN (n_29), .A (slo__sro_n321), .B1 (slo__sro_n322), .B2 (slo__sro_n320));
XNOR2_X1 slo__sro_c231 (.ZN (slo__sro_n319), .A (p_1[28]), .B (p_0[28]));
XNOR2_X1 slo__sro_c232 (.ZN (p_2[28]), .A (n_28), .B (slo__sro_n319));
OAI21_X1 slo__c248 (.ZN (slo__n339), .A (slo__sro_n65), .B1 (slo__sro_n66), .B2 (slo__sro_n64));
NAND2_X2 slo__sro_c363 (.ZN (n_22), .A1 (CLOCK_slo__sro_n1532), .A2 (slo__sro_n474));
XNOR2_X1 slo__sro_c364 (.ZN (slo__sro_n472), .A (p_1[21]), .B (p_0[21]));
XNOR2_X1 slo__sro_c365 (.ZN (p_2[21]), .A (slo__sro_n472), .B (n_21));
NOR2_X1 slo__sro_c374 (.ZN (slo__sro_n484), .A1 (n_33), .A2 (p_0[30]));
NAND2_X1 slo__sro_c375 (.ZN (slo__sro_n483), .A1 (slo__sro_n485), .A2 (slo__sro_n484));
OR2_X1 slo__sro_c376 (.ZN (slo__sro_n482), .A1 (p_1[30]), .A2 (n_34));
OAI21_X1 slo__sro_c377 (.ZN (slo__sro_n481), .A (slo__sro_n483), .B1 (n_32), .B2 (slo__sro_n482));
NAND2_X1 slo__sro_c437 (.ZN (slo__sro_n607), .A1 (p_1[5]), .A2 (p_0[5]));
NOR2_X1 slo__sro_c438 (.ZN (slo__sro_n606), .A1 (p_1[5]), .A2 (p_0[5]));
OAI21_X1 slo__sro_c439 (.ZN (slo__sro_n605), .A (slo__sro_n607), .B1 (slo__sro_n608), .B2 (slo__sro_n606));
NAND2_X1 CLOCK_slo__sro_c829 (.ZN (CLOCK_slo__sro_n1219), .A1 (p_1[2]), .A2 (p_0[2]));
NAND2_X1 slo__sro_c300 (.ZN (slo__sro_n405), .A1 (p_1[19]), .A2 (p_0[19]));
NOR2_X2 slo__sro_c301 (.ZN (slo__sro_n404), .A1 (p_1[19]), .A2 (p_0[19]));
OAI21_X1 slo__sro_c302 (.ZN (n_20), .A (slo__sro_n405), .B1 (slo__n869), .B2 (slo__sro_n404));
XNOR2_X1 slo__sro_c303 (.ZN (slo__sro_n403), .A (p_1[19]), .B (p_0[19]));
XNOR2_X1 slo__sro_c304 (.ZN (p_2[19]), .A (slo__sro_n171), .B (slo__sro_n403));
XNOR2_X1 slo__sro_c441 (.ZN (p_2[5]), .A (slo__sro_n604), .B (slo__sro_n216));
XNOR2_X1 slo__mro_c462 (.ZN (p_2[4]), .A (slo__mro_n638), .B (n_4));
INV_X1 CLOCK_slo__sro_c828 (.ZN (CLOCK_slo__sro_n1220), .A (n_2));
INV_X1 slo__L1_c630 (.ZN (slo__n869), .A (slo__sro_n171));
NOR2_X1 CLOCK_slo__sro_c830 (.ZN (CLOCK_slo__sro_n1218), .A1 (p_1[2]), .A2 (p_0[2]));
OAI21_X1 CLOCK_slo__sro_c831 (.ZN (CLOCK_slo__sro_n1217), .A (CLOCK_slo__sro_n1219)
    , .B1 (CLOCK_slo__sro_n1220), .B2 (CLOCK_slo__sro_n1218));
INV_X1 slo__sro_c713 (.ZN (slo__sro_n999), .A (n_22));
NAND2_X1 slo__sro_c714 (.ZN (slo__sro_n998), .A1 (p_1[22]), .A2 (p_0[22]));
NOR2_X1 slo__sro_c715 (.ZN (slo__sro_n997), .A1 (p_1[22]), .A2 (p_0[22]));
XNOR2_X1 slo__sro_c717 (.ZN (slo__sro_n996), .A (p_1[22]), .B (p_0[22]));
XNOR2_X1 slo__sro_c718 (.ZN (p_2[22]), .A (slo__sro_n996), .B (n_22));
XNOR2_X1 CLOCK_slo__sro_c833 (.ZN (p_2[2]), .A (n_2), .B (CLOCK_slo__sro_n1216));
NAND2_X1 CLOCK_slo__sro_c934 (.ZN (CLOCK_slo__sro_n1328), .A1 (p_1[15]), .A2 (p_0[15]));
NOR2_X1 CLOCK_slo__sro_c935 (.ZN (CLOCK_slo__sro_n1327), .A1 (p_1[15]), .A2 (p_0[15]));
OAI21_X2 CLOCK_slo__sro_c936 (.ZN (CLOCK_slo__sro_n1326), .A (CLOCK_slo__sro_n1328)
    , .B1 (CLOCK_slo__sro_n1329), .B2 (CLOCK_slo__sro_n1327));
XNOR2_X1 CLOCK_slo__sro_c937 (.ZN (CLOCK_slo__sro_n1325), .A (p_1[15]), .B (p_0[15]));
XNOR2_X1 CLOCK_slo__sro_c938 (.ZN (p_2[15]), .A (CLOCK_slo__sro_n1325), .B (n_15));
NAND2_X1 CLOCK_slo__sro_c1131 (.ZN (CLOCK_slo__sro_n1533), .A1 (CLOCK_slo__sro_n1535), .A2 (CLOCK_slo__sro_n1534));
OAI21_X2 CLOCK_slo__sro_c1066 (.ZN (n_12), .A (slo__sro_n204), .B1 (slo__sro_n205), .B2 (slo__sro_n203));
INV_X1 CLOCK_slo__sro_c1130 (.ZN (CLOCK_slo__sro_n1534), .A (p_0[21]));
NAND2_X1 CLOCK_slo__sro_c1132 (.ZN (CLOCK_slo__sro_n1532), .A1 (n_21), .A2 (CLOCK_slo__sro_n1533));
INV_X1 CLOCK_slo__sro_c986 (.ZN (CLOCK_slo__sro_n1388), .A (n_24));
NAND2_X1 CLOCK_slo__sro_c987 (.ZN (CLOCK_slo__sro_n1387), .A1 (p_1[24]), .A2 (p_0[24]));
NOR2_X1 CLOCK_slo__sro_c988 (.ZN (CLOCK_slo__sro_n1386), .A1 (p_1[24]), .A2 (p_0[24]));
OAI21_X1 CLOCK_slo__sro_c989 (.ZN (n_25), .A (CLOCK_slo__sro_n1387), .B1 (CLOCK_slo__sro_n1388), .B2 (CLOCK_slo__sro_n1386));
XNOR2_X1 CLOCK_slo__sro_c990 (.ZN (CLOCK_slo__sro_n1385), .A (p_1[24]), .B (p_0[24]));
XNOR2_X1 CLOCK_slo__sro_c991 (.ZN (p_2[24]), .A (CLOCK_slo__sro_n1385), .B (n_24));

endmodule //datapath__0_217

module datapath__0_216 (Multiplier_13_PP_0, Multiplier, p_0, p_1);

output [31:0] p_1;
input [31:0] Multiplier;
input [31:0] p_0;
input Multiplier_13_PP_0;
wire spw__n1757;
wire slo__sro_n550;
wire CLOCK_slo__sro_n1436;
wire slo__xsl_n773;
wire n_1;
wire n_2;
wire n_4;
wire n_6;
wire n_7;
wire n_8;
wire n_9;
wire n_10;
wire n_11;
wire n_12;
wire CLOCK_slo__sro_n1406;
wire n_16;
wire slo__sro_n498;
wire n_20;
wire n_21;
wire n_24;
wire n_26;
wire n_27;
wire n_30;
wire n_32;
wire n_0;
wire n_34;
wire n_33;
wire n_31;
wire slo__sro_n59;
wire slo__sro_n60;
wire slo__sro_n61;
wire slo__sro_n62;
wire slo__sro_n63;
wire slo__sro_n76;
wire slo__sro_n77;
wire slo__sro_n78;
wire slo__sro_n79;
wire slo__sro_n80;
wire slo__sro_n94;
wire slo__sro_n95;
wire slo__sro_n96;
wire slo__sro_n97;
wire slo__sro_n110;
wire slo__sro_n111;
wire slo__sro_n112;
wire slo__sro_n113;
wire slo__sro_n123;
wire slo__sro_n124;
wire slo__sro_n125;
wire slo__sro_n126;
wire slo__sro_n127;
wire slo__sro_n140;
wire slo__sro_n141;
wire slo__sro_n142;
wire slo__sro_n143;
wire slo__sro_n153;
wire slo__sro_n154;
wire slo__sro_n155;
wire slo__sro_n156;
wire slo__sro_n166;
wire slo__sro_n167;
wire slo__sro_n168;
wire slo__sro_n169;
wire slo__sro_n170;
wire slo__sro_n185;
wire slo__sro_n186;
wire slo__sro_n187;
wire slo__sro_n188;
wire slo__sro_n200;
wire slo__sro_n201;
wire slo__sro_n202;
wire slo__sro_n203;
wire slo__sro_n204;
wire slo__sro_n222;
wire slo__sro_n223;
wire slo__sro_n224;
wire slo__sro_n225;
wire slo__sro_n226;
wire slo__sro_n239;
wire slo__sro_n240;
wire slo__sro_n241;
wire slo__sro_n253;
wire slo__sro_n254;
wire slo__sro_n255;
wire slo__sro_n256;
wire slo__sro_n271;
wire slo__sro_n272;
wire slo__sro_n273;
wire slo__sro_n274;
wire slo__sro_n383;
wire slo__sro_n384;
wire slo__sro_n385;
wire slo__sro_n386;
wire slo__sro_n387;
wire slo__sro_n499;
wire slo__sro_n500;
wire slo__sro_n501;
wire slo__sro_n502;
wire slo__sro_n551;
wire slo__sro_n552;
wire slo__sro_n553;
wire slo__sro_n554;
wire slo__sro_n555;
wire slo__sro_n579;
wire slo__sro_n580;
wire slo__sro_n581;
wire slo__sro_n582;
wire slo__xsl_n774;
wire slo__sro_n1112;
wire slo__sro_n1113;
wire slo__sro_n1114;
wire slo__sro_n1115;
wire slo__sro_n1136;
wire slo__sro_n1137;
wire slo__sro_n1138;
wire slo__sro_n1139;
wire slo__sro_n1140;
wire CLOCK_slo__mro_n1391;
wire CLOCK_slo__sro_n1407;
wire CLOCK_slo__sro_n1408;
wire CLOCK_slo__sro_n1409;
wire CLOCK_slo__mro_n1423;
wire CLOCK_slo__sro_n1437;
wire CLOCK_slo__sro_n1438;
wire CLOCK_slo__sro_n1493;
wire CLOCK_slo__sro_n1494;
wire CLOCK_slo__sro_n1495;
wire CLOCK_slo__sro_n1496;


INV_X1 i_36 (.ZN (n_34), .A (Multiplier[30]));
INV_X1 i_35 (.ZN (n_33), .A (p_0[30]));
INV_X1 i_34 (.ZN (n_32), .A (n_30));
INV_X1 slo__sro_c745 (.ZN (slo__sro_n1140), .A (slo__sro_n124));
XOR2_X1 i_32 (.Z (p_1[31]), .A (Multiplier[31]), .B (n_31));
OAI22_X1 i_31 (.ZN (n_0), .A1 (n_34), .A2 (p_0[30]), .B1 (n_33), .B2 (Multiplier[30]));
XNOR2_X1 i_0 (.ZN (p_1[30]), .A (n_32), .B (n_0));
FA_X1 i_30 (.CO (n_30), .S (p_1[29]), .A (Multiplier[29]), .B (p_0[29]), .CI (slo__sro_n499));
INV_X1 slo__sro_c383 (.ZN (slo__sro_n554), .A (n_1));
INV_X1 slo__sro_c193 (.ZN (slo__sro_n274), .A (p_0[5]));
FA_X1 i_27 (.CO (n_27), .S (p_1[26]), .A (Multiplier[26]), .B (p_0[26]), .CI (n_26));
INV_X1 slo__sro_c177 (.ZN (slo__sro_n256), .A (n_27));
INV_X1 slo__sro_c115 (.ZN (slo__sro_n188), .A (n_9));
FA_X1 i_24 (.CO (n_24), .S (p_1[23]), .A (Multiplier[23]), .B (p_0[23]), .CI (slo__sro_n201));
INV_X1 slo__sro_c151 (.ZN (slo__sro_n226), .A (slo__sro_n384));
INV_X1 slo__xsl_c514 (.ZN (slo__xsl_n774), .A (slo__sro_n384));
INV_X1 slo__sro_c85 (.ZN (slo__sro_n156), .A (n_7));
XNOR2_X1 CLOCK_slo__mro_c928 (.ZN (CLOCK_slo__mro_n1423), .A (p_0[27]), .B (Multiplier[27]));
NAND2_X1 slo__sro_c165 (.ZN (slo__sro_n241), .A1 (slo__sro_n167), .A2 (Multiplier[25]));
NAND2_X1 slo__sro_c355 (.ZN (slo__sro_n501), .A1 (p_0[28]), .A2 (Multiplier[28]));
INV_X1 slo__sro_c15 (.ZN (slo__sro_n80), .A (slo__sro_n1137));
FA_X1 i_16 (.CO (n_16), .S (p_1[15]), .A (Multiplier[15]), .B (p_0[15]), .CI (slo__sro_n77));
INV_X1 slo__sro_c29 (.ZN (slo__sro_n97), .A (n_4));
CLKBUF_X2 spw__c1305 (.Z (slo__sro_n224), .A (spw__n1757));
INV_X2 slo__sro_c71 (.ZN (slo__sro_n143), .A (n_20));
FA_X1 i_12 (.CO (n_12), .S (p_1[11]), .A (Multiplier[11]), .B (p_0[11]), .CI (n_11));
INV_X1 slo__sro_c57 (.ZN (slo__sro_n127), .A (n_12));
INV_X1 slo__sro_c129 (.ZN (slo__sro_n204), .A (slo__sro_n580));
FA_X1 i_9 (.CO (n_9), .S (p_1[8]), .A (Multiplier[8]), .B (p_0[8]), .CI (n_8));
INV_X1 slo__sro_c99 (.ZN (slo__sro_n170), .A (n_24));
FA_X1 i_7 (.CO (n_7), .S (p_1[6]), .A (Multiplier[6]), .B (p_0[6]), .CI (n_6));
INV_X1 slo__sro_c382 (.ZN (slo__sro_n555), .A (Multiplier[1]));
INV_X1 slo__sro_c43 (.ZN (slo__sro_n113), .A (n_10));
NAND2_X1 CLOCK_slo__sro_c998 (.ZN (CLOCK_slo__sro_n1496), .A1 (p_0[2]), .A2 (Multiplier[2]));
NAND2_X1 slo__sro_c410 (.ZN (slo__sro_n582), .A1 (p_0[21]), .A2 (Multiplier[21]));
HA_X1 i_1 (.CO (n_1), .S (p_1[0]), .A (Multiplier[0]), .B (p_0[0]));
INV_X1 slo__sro_c1 (.ZN (slo__sro_n63), .A (n_16));
NAND2_X1 slo__sro_c2 (.ZN (slo__sro_n62), .A1 (p_0[16]), .A2 (Multiplier[16]));
NOR2_X1 slo__sro_c3 (.ZN (slo__sro_n61), .A1 (p_0[16]), .A2 (Multiplier[16]));
OAI21_X2 slo__sro_c4 (.ZN (slo__sro_n60), .A (slo__sro_n62), .B1 (slo__sro_n61), .B2 (slo__sro_n63));
XNOR2_X2 slo__sro_c5 (.ZN (slo__sro_n59), .A (p_0[16]), .B (Multiplier[16]));
XNOR2_X1 slo__sro_c6 (.ZN (p_1[16]), .A (slo__sro_n59), .B (n_16));
NAND2_X1 slo__sro_c16 (.ZN (slo__sro_n79), .A1 (p_0[14]), .A2 (Multiplier[14]));
NOR2_X1 slo__sro_c17 (.ZN (slo__sro_n78), .A1 (p_0[14]), .A2 (Multiplier[14]));
OAI21_X1 slo__sro_c18 (.ZN (slo__sro_n77), .A (slo__sro_n79), .B1 (slo__sro_n80), .B2 (slo__sro_n78));
XNOR2_X1 slo__sro_c19 (.ZN (slo__sro_n76), .A (p_0[14]), .B (Multiplier[14]));
XNOR2_X1 slo__sro_c20 (.ZN (p_1[14]), .A (slo__sro_n76), .B (slo__sro_n1137));
NAND2_X1 slo__sro_c30 (.ZN (slo__sro_n96), .A1 (p_0[4]), .A2 (Multiplier[4]));
NOR2_X1 slo__sro_c31 (.ZN (slo__sro_n95), .A1 (p_0[4]), .A2 (Multiplier[4]));
OAI21_X2 slo__sro_c32 (.ZN (slo__sro_n94), .A (slo__sro_n96), .B1 (slo__sro_n95), .B2 (slo__sro_n97));
INV_X2 CLOCK_slo__sro_c909 (.ZN (CLOCK_slo__sro_n1409), .A (slo__sro_n223));
NAND2_X1 CLOCK_slo__sro_c910 (.ZN (CLOCK_slo__sro_n1408), .A1 (p_0[19]), .A2 (Multiplier[19]));
NAND2_X1 slo__sro_c44 (.ZN (slo__sro_n112), .A1 (p_0[10]), .A2 (Multiplier[10]));
NOR2_X1 slo__sro_c45 (.ZN (slo__sro_n111), .A1 (p_0[10]), .A2 (Multiplier[10]));
OAI21_X1 slo__sro_c46 (.ZN (n_11), .A (slo__sro_n112), .B1 (slo__sro_n111), .B2 (slo__sro_n113));
XNOR2_X1 slo__sro_c47 (.ZN (slo__sro_n110), .A (p_0[10]), .B (Multiplier[10]));
XNOR2_X1 slo__sro_c48 (.ZN (p_1[10]), .A (slo__sro_n110), .B (n_10));
NAND2_X1 slo__sro_c58 (.ZN (slo__sro_n126), .A1 (p_0[12]), .A2 (Multiplier[12]));
NOR2_X1 slo__sro_c59 (.ZN (slo__sro_n125), .A1 (p_0[12]), .A2 (Multiplier[12]));
OAI21_X1 slo__sro_c60 (.ZN (slo__sro_n124), .A (slo__sro_n126), .B1 (slo__sro_n127), .B2 (slo__sro_n125));
XNOR2_X2 slo__sro_c61 (.ZN (slo__sro_n123), .A (p_0[12]), .B (Multiplier[12]));
XNOR2_X1 slo__sro_c62 (.ZN (p_1[12]), .A (slo__sro_n123), .B (n_12));
NAND2_X1 slo__sro_c72 (.ZN (slo__sro_n142), .A1 (p_0[20]), .A2 (Multiplier[20]));
NOR2_X1 slo__sro_c73 (.ZN (slo__sro_n141), .A1 (p_0[20]), .A2 (Multiplier[20]));
OAI21_X2 slo__sro_c74 (.ZN (n_21), .A (slo__sro_n142), .B1 (slo__sro_n143), .B2 (slo__sro_n141));
XNOR2_X1 slo__sro_c75 (.ZN (slo__sro_n140), .A (p_0[20]), .B (Multiplier[20]));
XNOR2_X1 slo__sro_c76 (.ZN (p_1[20]), .A (slo__sro_n140), .B (n_20));
NAND2_X1 slo__sro_c86 (.ZN (slo__sro_n155), .A1 (p_0[7]), .A2 (Multiplier[7]));
NOR2_X1 slo__sro_c87 (.ZN (slo__sro_n154), .A1 (p_0[7]), .A2 (Multiplier[7]));
OAI21_X1 slo__sro_c88 (.ZN (n_8), .A (slo__sro_n155), .B1 (slo__sro_n156), .B2 (slo__sro_n154));
XNOR2_X1 slo__sro_c89 (.ZN (slo__sro_n153), .A (p_0[7]), .B (Multiplier[7]));
XNOR2_X1 slo__sro_c90 (.ZN (p_1[7]), .A (slo__sro_n153), .B (n_7));
NAND2_X1 slo__sro_c100 (.ZN (slo__sro_n169), .A1 (p_0[24]), .A2 (Multiplier[24]));
NOR2_X1 slo__sro_c101 (.ZN (slo__sro_n168), .A1 (p_0[24]), .A2 (Multiplier[24]));
OAI21_X2 slo__sro_c102 (.ZN (slo__sro_n167), .A (slo__sro_n169), .B1 (slo__sro_n170), .B2 (slo__sro_n168));
XNOR2_X2 slo__sro_c103 (.ZN (slo__sro_n166), .A (p_0[24]), .B (Multiplier[24]));
XNOR2_X1 slo__sro_c104 (.ZN (p_1[24]), .A (slo__sro_n166), .B (n_24));
NAND2_X1 slo__sro_c116 (.ZN (slo__sro_n187), .A1 (p_0[9]), .A2 (Multiplier[9]));
NOR2_X1 slo__sro_c117 (.ZN (slo__sro_n186), .A1 (p_0[9]), .A2 (Multiplier[9]));
OAI21_X1 slo__sro_c118 (.ZN (n_10), .A (slo__sro_n187), .B1 (slo__sro_n188), .B2 (slo__sro_n186));
XNOR2_X1 slo__sro_c119 (.ZN (slo__sro_n185), .A (p_0[9]), .B (Multiplier[9]));
XNOR2_X1 slo__sro_c120 (.ZN (p_1[9]), .A (slo__sro_n185), .B (n_9));
NAND2_X1 slo__sro_c130 (.ZN (slo__sro_n203), .A1 (p_0[22]), .A2 (Multiplier[22]));
NOR2_X2 slo__sro_c131 (.ZN (slo__sro_n202), .A1 (p_0[22]), .A2 (Multiplier[22]));
OAI21_X1 slo__sro_c132 (.ZN (slo__sro_n201), .A (slo__sro_n203), .B1 (slo__sro_n202), .B2 (slo__sro_n204));
XNOR2_X1 slo__sro_c133 (.ZN (slo__sro_n200), .A (p_0[22]), .B (Multiplier[22]));
XNOR2_X1 slo__sro_c134 (.ZN (p_1[22]), .A (slo__sro_n200), .B (slo__sro_n580));
NAND2_X1 slo__sro_c152 (.ZN (slo__sro_n225), .A1 (p_0[18]), .A2 (Multiplier[18]));
NOR2_X1 slo__sro_c153 (.ZN (spw__n1757), .A1 (p_0[18]), .A2 (Multiplier[18]));
INV_X1 slo__sro_c719 (.ZN (slo__sro_n1115), .A (n_30));
XNOR2_X2 slo__sro_c155 (.ZN (slo__sro_n222), .A (p_0[18]), .B (Multiplier[18]));
XNOR2_X2 slo__sro_c156 (.ZN (p_1[18]), .A (slo__sro_n222), .B (slo__xsl_n773));
OAI21_X1 slo__sro_c166 (.ZN (slo__sro_n240), .A (p_0[25]), .B1 (slo__sro_n167), .B2 (Multiplier[25]));
NAND2_X1 slo__sro_c167 (.ZN (n_26), .A1 (slo__sro_n240), .A2 (slo__sro_n241));
XNOR2_X2 slo__sro_c168 (.ZN (slo__sro_n239), .A (slo__sro_n167), .B (Multiplier[25]));
XNOR2_X2 slo__sro_c169 (.ZN (p_1[25]), .A (slo__sro_n239), .B (p_0[25]));
NAND2_X1 slo__sro_c178 (.ZN (slo__sro_n255), .A1 (p_0[27]), .A2 (Multiplier[27]));
NOR2_X1 slo__sro_c179 (.ZN (slo__sro_n254), .A1 (p_0[27]), .A2 (Multiplier[27]));
OAI21_X4 slo__sro_c180 (.ZN (slo__sro_n253), .A (slo__sro_n255), .B1 (slo__sro_n254), .B2 (slo__sro_n256));
NAND2_X1 CLOCK_slo__sro_c938 (.ZN (CLOCK_slo__sro_n1438), .A1 (p_0[3]), .A2 (Multiplier[3]));
OAI21_X2 CLOCK_slo__sro_c939 (.ZN (CLOCK_slo__sro_n1437), .A (CLOCK_slo__sro_n1494)
    , .B1 (p_0[3]), .B2 (Multiplier[3]));
NAND2_X1 slo__sro_c194 (.ZN (slo__sro_n273), .A1 (slo__sro_n94), .A2 (Multiplier[5]));
NOR2_X1 slo__sro_c195 (.ZN (slo__sro_n272), .A1 (slo__sro_n94), .A2 (Multiplier[5]));
OAI21_X1 slo__sro_c196 (.ZN (n_6), .A (slo__sro_n273), .B1 (slo__sro_n272), .B2 (slo__sro_n274));
XNOR2_X1 slo__sro_c197 (.ZN (slo__sro_n271), .A (slo__sro_n94), .B (Multiplier[5]));
XNOR2_X1 slo__sro_c198 (.ZN (p_1[5]), .A (slo__sro_n271), .B (p_0[5]));
INV_X1 slo__sro_c354 (.ZN (slo__sro_n502), .A (slo__sro_n253));
INV_X1 slo__sro_c266 (.ZN (slo__sro_n387), .A (slo__sro_n60));
NAND2_X1 slo__sro_c267 (.ZN (slo__sro_n386), .A1 (p_0[17]), .A2 (Multiplier[17]));
NOR2_X2 slo__sro_c268 (.ZN (slo__sro_n385), .A1 (p_0[17]), .A2 (Multiplier[17]));
OAI21_X2 slo__sro_c269 (.ZN (slo__sro_n384), .A (slo__sro_n386), .B1 (slo__sro_n387), .B2 (slo__sro_n385));
XNOR2_X2 slo__sro_c270 (.ZN (slo__sro_n383), .A (p_0[17]), .B (Multiplier[17]));
XNOR2_X1 slo__sro_c271 (.ZN (p_1[17]), .A (slo__sro_n383), .B (slo__sro_n60));
NOR2_X1 slo__sro_c356 (.ZN (slo__sro_n500), .A1 (p_0[28]), .A2 (Multiplier[28]));
OAI21_X2 slo__sro_c357 (.ZN (slo__sro_n499), .A (slo__sro_n501), .B1 (slo__sro_n502), .B2 (slo__sro_n500));
XNOR2_X1 slo__sro_c358 (.ZN (slo__sro_n498), .A (p_0[28]), .B (Multiplier[28]));
XNOR2_X1 slo__sro_c359 (.ZN (p_1[28]), .A (slo__sro_n498), .B (slo__sro_n253));
NAND2_X1 slo__sro_c384 (.ZN (slo__sro_n553), .A1 (n_1), .A2 (Multiplier[1]));
NAND2_X1 slo__sro_c385 (.ZN (slo__sro_n552), .A1 (slo__sro_n554), .A2 (slo__sro_n555));
NAND2_X1 slo__sro_c386 (.ZN (slo__sro_n551), .A1 (p_0[1]), .A2 (slo__sro_n552));
NAND2_X1 slo__sro_c387 (.ZN (n_2), .A1 (slo__sro_n551), .A2 (slo__sro_n553));
XNOR2_X1 slo__sro_c388 (.ZN (slo__sro_n550), .A (n_1), .B (Multiplier[1]));
XNOR2_X1 slo__sro_c389 (.ZN (p_1[1]), .A (p_0[1]), .B (slo__sro_n550));
OAI21_X1 slo__sro_c411 (.ZN (slo__sro_n581), .A (n_21), .B1 (p_0[21]), .B2 (Multiplier[21]));
NAND2_X2 slo__sro_c412 (.ZN (slo__sro_n580), .A1 (slo__sro_n581), .A2 (slo__sro_n582));
XNOR2_X2 slo__sro_c413 (.ZN (slo__sro_n579), .A (n_21), .B (Multiplier[21]));
XNOR2_X1 slo__sro_c414 (.ZN (p_1[21]), .A (slo__sro_n579), .B (p_0[21]));
INV_X1 slo__xsl_c515 (.ZN (slo__xsl_n773), .A (slo__xsl_n774));
OAI21_X4 slo__sro_c695 (.ZN (slo__sro_n223), .A (slo__sro_n225), .B1 (slo__sro_n226), .B2 (slo__sro_n224));
NOR2_X1 slo__sro_c720 (.ZN (slo__sro_n1114), .A1 (n_33), .A2 (Multiplier[30]));
NAND2_X1 slo__sro_c721 (.ZN (slo__sro_n1113), .A1 (slo__sro_n1114), .A2 (slo__sro_n1115));
OR2_X1 slo__sro_c722 (.ZN (slo__sro_n1112), .A1 (p_0[30]), .A2 (n_34));
OAI21_X1 slo__sro_c723 (.ZN (n_31), .A (slo__sro_n1113), .B1 (n_32), .B2 (slo__sro_n1112));
NAND2_X1 slo__sro_c746 (.ZN (slo__sro_n1139), .A1 (p_0[13]), .A2 (Multiplier[13]));
NOR2_X2 slo__sro_c747 (.ZN (slo__sro_n1138), .A1 (p_0[13]), .A2 (Multiplier_13_PP_0));
OAI21_X2 slo__sro_c748 (.ZN (slo__sro_n1137), .A (slo__sro_n1139), .B1 (slo__sro_n1140), .B2 (slo__sro_n1138));
XNOR2_X1 slo__sro_c749 (.ZN (slo__sro_n1136), .A (p_0[13]), .B (Multiplier[13]));
XNOR2_X1 slo__sro_c750 (.ZN (p_1[13]), .A (slo__sro_n1136), .B (slo__sro_n124));
XNOR2_X1 CLOCK_slo__mro_c897 (.ZN (CLOCK_slo__mro_n1391), .A (n_4), .B (Multiplier[4]));
XNOR2_X1 CLOCK_slo__mro_c898 (.ZN (p_1[4]), .A (CLOCK_slo__mro_n1391), .B (p_0[4]));
NOR2_X1 CLOCK_slo__sro_c911 (.ZN (CLOCK_slo__sro_n1407), .A1 (p_0[19]), .A2 (Multiplier[19]));
OAI21_X2 CLOCK_slo__sro_c912 (.ZN (n_20), .A (CLOCK_slo__sro_n1408), .B1 (CLOCK_slo__sro_n1407), .B2 (CLOCK_slo__sro_n1409));
XNOR2_X2 CLOCK_slo__sro_c913 (.ZN (CLOCK_slo__sro_n1406), .A (p_0[19]), .B (Multiplier[19]));
XNOR2_X2 CLOCK_slo__sro_c914 (.ZN (p_1[19]), .A (CLOCK_slo__sro_n1406), .B (slo__sro_n223));
XNOR2_X1 CLOCK_slo__mro_c929 (.ZN (p_1[27]), .A (CLOCK_slo__mro_n1423), .B (n_27));
NAND2_X2 CLOCK_slo__sro_c940 (.ZN (n_4), .A1 (CLOCK_slo__sro_n1437), .A2 (CLOCK_slo__sro_n1438));
XNOR2_X1 CLOCK_slo__sro_c941 (.ZN (CLOCK_slo__sro_n1436), .A (CLOCK_slo__sro_n1494), .B (Multiplier[3]));
XNOR2_X1 CLOCK_slo__sro_c942 (.ZN (p_1[3]), .A (CLOCK_slo__sro_n1436), .B (p_0[3]));
OAI21_X2 CLOCK_slo__sro_c999 (.ZN (CLOCK_slo__sro_n1495), .A (n_2), .B1 (p_0[2]), .B2 (Multiplier[2]));
NAND2_X4 CLOCK_slo__sro_c1000 (.ZN (CLOCK_slo__sro_n1494), .A1 (CLOCK_slo__sro_n1495), .A2 (CLOCK_slo__sro_n1496));
XNOR2_X2 CLOCK_slo__sro_c1001 (.ZN (CLOCK_slo__sro_n1493), .A (p_0[2]), .B (Multiplier[2]));
XNOR2_X2 CLOCK_slo__sro_c1002 (.ZN (p_1[2]), .A (CLOCK_slo__sro_n1493), .B (n_2));

endmodule //datapath__0_216

module datapath__0_212 (opt_ipoPP_2, p_0, p_1, p_2);

output [31:0] p_2;
input [31:0] p_0;
input [31:0] p_1;
input opt_ipoPP_2;
wire slo__sro_n941;
wire n_1;
wire slo__sro_n1024;
wire n_3;
wire n_4;
wire n_5;
wire n_6;
wire n_7;
wire n_8;
wire n_9;
wire n_10;
wire n_11;
wire n_12;
wire slo__sro_n355;
wire n_14;
wire n_15;
wire CLOCK_slo__sro_n1531;
wire n_17;
wire n_18;
wire n_20;
wire n_21;
wire n_23;
wire n_24;
wire n_26;
wire n_27;
wire n_28;
wire n_29;
wire n_30;
wire n_32;
wire n_0;
wire n_34;
wire n_33;
wire n_31;
wire slo__sro_n65;
wire slo__sro_n66;
wire slo__sro_n67;
wire slo__sro_n68;
wire slo__sro_n338;
wire slo__sro_n339;
wire slo__sro_n340;
wire slo__sro_n341;
wire slo__sro_n342;
wire CLOCK_slo__sro_n1430;
wire slo__sro_n321;
wire slo__sro_n322;
wire slo__sro_n323;
wire slo__sro_n324;
wire slo__sro_n325;
wire slo__sro_n356;
wire slo__sro_n357;
wire slo__sro_n358;
wire slo__sro_n380;
wire slo__sro_n381;
wire slo__sro_n383;
wire slo__sro_n435;
wire slo__sro_n436;
wire slo__sro_n437;
wire slo__sro_n438;
wire slo__sro_n598;
wire slo__sro_n599;
wire slo__sro_n600;
wire slo__sro_n601;
wire slo__sro_n942;
wire slo__sro_n943;
wire slo__sro_n944;
wire slo__sro_n1020;
wire slo__sro_n1021;
wire slo__sro_n1022;
wire slo__sro_n1023;
wire slo__sro_n667;
wire slo__sro_n668;
wire slo__sro_n669;
wire slo__sro_n670;
wire CLOCK_slo__sro_n1431;
wire CLOCK_slo__sro_n1432;
wire CLOCK_slo__sro_n1433;
wire CLOCK_slo__sro_n1434;
wire CLOCK_slo__mro_n1886;
wire slo__sro_n1099;
wire slo__sro_n1100;
wire slo__sro_n1101;
wire slo__sro_n1102;
wire CLOCK_slo__sro_n1529;
wire CLOCK_slo__sro_n1530;
wire CLOCK_slo__sro_n1467;
wire CLOCK_slo__sro_n1468;
wire CLOCK_slo__sro_n1470;
wire CLOCK_slo__sro_n1471;
wire CLOCK_slo__sro_n1548;
wire CLOCK_slo__sro_n1549;
wire CLOCK_slo__sro_n1550;
wire CLOCK_slo__sro_n1551;
wire CLOCK_slo__sro_n1559;
wire CLOCK_slo__sro_n1633;
wire CLOCK_slo__sro_n1634;
wire CLOCK_slo__sro_n1635;
wire CLOCK_slo__sro_n1592;
wire CLOCK_slo__sro_n1593;
wire CLOCK_slo__sro_n1594;
wire CLOCK_slo__sro_n1806;
wire CLOCK_slo__sro_n1805;
wire CLOCK_slo__sro_n1807;
wire CLOCK_slo__sro_n1808;


INV_X1 i_36 (.ZN (n_34), .A (p_0[30]));
INV_X1 i_35 (.ZN (n_33), .A (p_1[30]));
INV_X1 i_34 (.ZN (n_32), .A (n_30));
XOR2_X1 i_32 (.Z (p_2[31]), .A (n_31), .B (p_0[31]));
OAI22_X1 i_31 (.ZN (n_0), .A1 (n_34), .A2 (p_1[30]), .B1 (p_0[30]), .B2 (n_33));
XNOR2_X1 i_0 (.ZN (p_2[30]), .A (n_32), .B (n_0));
NAND2_X1 slo__sro_c698 (.ZN (slo__sro_n943), .A1 (p_1[7]), .A2 (p_0[7]));
FA_X1 i_29 (.CO (n_29), .S (p_2[28]), .A (p_0[28]), .B (p_1[28]), .CI (n_28));
INV_X1 CLOCK_slo__sro_c1112 (.ZN (CLOCK_slo__sro_n1551), .A (n_6));
FA_X1 i_27 (.CO (n_27), .S (p_2[26]), .A (p_0[26]), .B (p_1[26]), .CI (n_26));
FA_X1 i_26 (.CO (n_26), .S (p_2[25]), .A (p_0[25]), .B (p_1[25]), .CI (slo__sro_n381));
INV_X1 slo__sro_c359 (.ZN (slo__sro_n438), .A (n_8));
INV_X1 slo__sro_c267 (.ZN (slo__sro_n342), .A (n_18));
FA_X1 i_23 (.CO (n_23), .S (p_2[22]), .A (p_0[22]), .B (p_1[22]), .CI (slo__sro_n1021));
XNOR2_X2 slo__sro_c885 (.ZN (p_2[12]), .A (slo__sro_n321), .B (n_12));
FA_X1 i_21 (.CO (n_21), .S (p_2[20]), .A (p_0[20]), .B (p_1[20]), .CI (n_20));
NAND2_X1 slo__sro_c308 (.ZN (slo__sro_n383), .A1 (p_1[24]), .A2 (p_0[24]));
INV_X1 slo__sro_c281 (.ZN (slo__sro_n358), .A (slo__sro_n339));
NAND2_X1 CLOCK_slo__sro_c1093 (.ZN (n_28), .A1 (CLOCK_slo__sro_n1530), .A2 (CLOCK_slo__sro_n1531));
XNOR2_X1 CLOCK_slo__sro_c1095 (.ZN (p_2[27]), .A (CLOCK_slo__sro_n1529), .B (n_27));
FA_X1 i_15 (.CO (n_15), .S (p_2[14]), .A (p_0[14]), .B (p_1[14]), .CI (n_14));
FA_X1 i_14 (.CO (n_14), .S (p_2[13]), .A (p_0[13]), .B (p_1[13]), .CI (slo__sro_n322));
NAND2_X1 slo__sro_c282 (.ZN (slo__sro_n357), .A1 (p_1[19]), .A2 (p_0[19]));
FA_X1 i_12 (.CO (n_12), .S (p_2[11]), .A (p_0[11]), .B (p_1[11]), .CI (n_11));
INV_X1 CLOCK_slo__sro_c1347 (.ZN (CLOCK_slo__sro_n1808), .A (n_17));
INV_X1 slo__sro_c697 (.ZN (slo__sro_n944), .A (n_7));
INV_X1 slo__sro_c772 (.ZN (slo__sro_n1024), .A (n_21));
OAI21_X1 CLOCK_slo__sro_c1126 (.ZN (CLOCK_slo__sro_n1559), .A (n_24), .B1 (p_1[24]), .B2 (p_0[24]));
FA_X1 i_6 (.CO (n_6), .S (p_2[5]), .A (p_0[5]), .B (p_1[5]), .CI (n_5));
FA_X1 i_5 (.CO (n_5), .S (p_2[4]), .A (p_0[4]), .B (p_1[4]), .CI (n_4));
FA_X1 i_4 (.CO (n_4), .S (p_2[3]), .A (p_0[3]), .B (p_1[3]), .CI (n_3));
FA_X1 i_3 (.CO (n_3), .S (p_2[2]), .A (p_0[2]), .B (p_1[2]), .CI (slo__sro_n668));
NOR2_X1 CLOCK_slo__sro_c991 (.ZN (CLOCK_slo__sro_n1431), .A1 (p_1[30]), .A2 (n_34));
HA_X1 i_1 (.CO (n_1), .S (p_2[0]), .A (p_0[0]), .B (p_1[0]));
INV_X1 slo__sro_c3 (.ZN (slo__sro_n68), .A (n_23));
NAND2_X1 slo__sro_c4 (.ZN (slo__sro_n67), .A1 (p_1[23]), .A2 (p_0[23]));
NOR2_X1 slo__sro_c5 (.ZN (slo__sro_n66), .A1 (p_1[23]), .A2 (p_0[23]));
OAI21_X2 slo__sro_c6 (.ZN (n_24), .A (slo__sro_n67), .B1 (slo__sro_n68), .B2 (slo__sro_n66));
XNOR2_X1 slo__sro_c7 (.ZN (slo__sro_n65), .A (p_1[23]), .B (p_0[23]));
XNOR2_X1 slo__sro_c8 (.ZN (p_2[23]), .A (slo__sro_n65), .B (n_23));
NAND2_X1 slo__sro_c268 (.ZN (slo__sro_n341), .A1 (p_1[18]), .A2 (p_0[18]));
NOR2_X1 slo__sro_c269 (.ZN (slo__sro_n340), .A1 (p_1[18]), .A2 (p_0[18]));
OAI21_X1 slo__sro_c270 (.ZN (slo__sro_n339), .A (slo__sro_n341), .B1 (slo__sro_n342), .B2 (slo__sro_n340));
XNOR2_X1 slo__sro_c271 (.ZN (slo__sro_n338), .A (p_1[18]), .B (p_0[18]));
XNOR2_X1 slo__sro_c272 (.ZN (p_2[18]), .A (slo__sro_n338), .B (n_18));
INV_X1 slo__sro_c253 (.ZN (slo__sro_n325), .A (n_12));
NAND2_X1 slo__sro_c254 (.ZN (slo__sro_n324), .A1 (p_1[12]), .A2 (p_0[12]));
NOR2_X1 slo__sro_c255 (.ZN (slo__sro_n323), .A1 (p_1[12]), .A2 (p_0[12]));
OAI21_X1 slo__sro_c256 (.ZN (slo__sro_n322), .A (slo__sro_n324), .B1 (slo__sro_n325), .B2 (slo__sro_n323));
XNOR2_X2 slo__sro_c257 (.ZN (slo__sro_n321), .A (p_1[12]), .B (p_0[12]));
NOR2_X1 CLOCK_slo__sro_c989 (.ZN (CLOCK_slo__sro_n1433), .A1 (n_30), .A2 (n_33));
NOR2_X1 slo__sro_c283 (.ZN (slo__sro_n356), .A1 (p_1[19]), .A2 (p_0[19]));
OAI21_X1 slo__sro_c284 (.ZN (n_20), .A (slo__sro_n357), .B1 (slo__sro_n358), .B2 (slo__sro_n356));
XNOR2_X1 slo__sro_c285 (.ZN (slo__sro_n355), .A (p_1[19]), .B (p_0[19]));
XNOR2_X1 slo__sro_c286 (.ZN (p_2[19]), .A (slo__sro_n355), .B (slo__sro_n339));
NOR2_X1 CLOCK_slo__mro_c1436 (.ZN (CLOCK_slo__mro_n1886), .A1 (p_1[15]), .A2 (p_0[15]));
NAND2_X1 slo__sro_c310 (.ZN (slo__sro_n381), .A1 (CLOCK_slo__sro_n1559), .A2 (slo__sro_n383));
XNOR2_X2 slo__sro_c311 (.ZN (slo__sro_n380), .A (n_24), .B (p_0[24]));
XNOR2_X2 slo__sro_c312 (.ZN (p_2[24]), .A (slo__sro_n380), .B (p_1[24]));
NAND2_X1 slo__sro_c360 (.ZN (slo__sro_n437), .A1 (p_1[8]), .A2 (p_0[8]));
NOR2_X1 slo__sro_c361 (.ZN (slo__sro_n436), .A1 (p_1[8]), .A2 (p_0[8]));
OAI21_X1 slo__sro_c362 (.ZN (n_9), .A (slo__sro_n437), .B1 (slo__sro_n436), .B2 (slo__sro_n438));
XNOR2_X2 slo__sro_c363 (.ZN (slo__sro_n435), .A (p_1[8]), .B (p_0[8]));
XNOR2_X1 slo__sro_c364 (.ZN (p_2[8]), .A (slo__sro_n435), .B (n_8));
INV_X1 slo__sro_c449 (.ZN (slo__sro_n601), .A (n_29));
NAND2_X1 slo__sro_c450 (.ZN (slo__sro_n600), .A1 (p_1[29]), .A2 (p_0[29]));
NOR2_X1 slo__sro_c451 (.ZN (slo__sro_n599), .A1 (p_1[29]), .A2 (p_0[29]));
NAND2_X1 CLOCK_slo__sro_c1348 (.ZN (CLOCK_slo__sro_n1807), .A1 (p_1[17]), .A2 (p_0[17]));
XNOR2_X1 slo__sro_c453 (.ZN (slo__sro_n598), .A (p_1[29]), .B (p_0[29]));
XNOR2_X1 slo__sro_c454 (.ZN (p_2[29]), .A (slo__sro_n598), .B (n_29));
NOR2_X1 slo__sro_c699 (.ZN (slo__sro_n942), .A1 (p_1[7]), .A2 (p_0[7]));
OAI21_X2 slo__sro_c700 (.ZN (n_8), .A (slo__sro_n943), .B1 (slo__sro_n944), .B2 (slo__sro_n942));
XNOR2_X1 slo__sro_c701 (.ZN (slo__sro_n941), .A (p_1[7]), .B (p_0[7]));
XNOR2_X1 slo__sro_c702 (.ZN (p_2[7]), .A (slo__sro_n941), .B (n_7));
NAND2_X1 slo__sro_c773 (.ZN (slo__sro_n1023), .A1 (p_1[21]), .A2 (p_0[21]));
NOR2_X1 slo__sro_c774 (.ZN (slo__sro_n1022), .A1 (p_1[21]), .A2 (p_0[21]));
OAI21_X1 slo__sro_c775 (.ZN (slo__sro_n1021), .A (slo__sro_n1023), .B1 (slo__sro_n1024), .B2 (slo__sro_n1022));
XNOR2_X1 slo__sro_c776 (.ZN (slo__sro_n1020), .A (p_1[21]), .B (p_0[21]));
XNOR2_X1 slo__sro_c777 (.ZN (p_2[21]), .A (slo__sro_n1020), .B (n_21));
NAND2_X1 CLOCK_slo__sro_c990 (.ZN (CLOCK_slo__sro_n1432), .A1 (CLOCK_slo__sro_n1433), .A2 (CLOCK_slo__sro_n1434));
INV_X1 CLOCK_slo__sro_c988 (.ZN (CLOCK_slo__sro_n1434), .A (p_0[30]));
NAND2_X1 slo__sro_c510 (.ZN (slo__sro_n670), .A1 (n_1), .A2 (p_0[1]));
NOR2_X1 slo__sro_c511 (.ZN (slo__sro_n669), .A1 (n_1), .A2 (p_0[1]));
OAI21_X1 slo__sro_c512 (.ZN (slo__sro_n668), .A (slo__sro_n670), .B1 (p_1[1]), .B2 (slo__sro_n669));
XNOR2_X1 slo__sro_c513 (.ZN (slo__sro_n667), .A (n_1), .B (p_0[1]));
XNOR2_X1 slo__sro_c514 (.ZN (p_2[1]), .A (opt_ipoPP_2), .B (slo__sro_n667));
INV_X1 CLOCK_slo__sro_c992 (.ZN (CLOCK_slo__sro_n1430), .A (CLOCK_slo__sro_n1431));
OAI21_X1 CLOCK_slo__sro_c993 (.ZN (n_31), .A (CLOCK_slo__sro_n1432), .B1 (n_32), .B2 (CLOCK_slo__sro_n1430));
NAND2_X1 CLOCK_slo__sro_c1091 (.ZN (CLOCK_slo__sro_n1531), .A1 (p_0[27]), .A2 (p_1[27]));
OAI21_X1 CLOCK_slo__sro_c1092 (.ZN (CLOCK_slo__sro_n1530), .A (n_27), .B1 (p_1[27]), .B2 (p_0[27]));
INV_X1 slo__sro_c839 (.ZN (slo__sro_n1102), .A (CLOCK_slo__sro_n1468));
NAND2_X1 slo__sro_c840 (.ZN (slo__sro_n1101), .A1 (p_1[16]), .A2 (p_0[16]));
NOR2_X1 slo__sro_c841 (.ZN (slo__sro_n1100), .A1 (p_1[16]), .A2 (p_0[16]));
OAI21_X1 slo__sro_c842 (.ZN (n_17), .A (slo__sro_n1101), .B1 (slo__sro_n1102), .B2 (slo__sro_n1100));
XNOR2_X1 slo__sro_c843 (.ZN (slo__sro_n1099), .A (p_1[16]), .B (p_0[16]));
XNOR2_X1 slo__sro_c844 (.ZN (p_2[16]), .A (slo__sro_n1099), .B (CLOCK_slo__sro_n1468));
XNOR2_X1 CLOCK_slo__sro_c1094 (.ZN (CLOCK_slo__sro_n1529), .A (p_1[27]), .B (p_0[27]));
INV_X1 CLOCK_slo__sro_c1028 (.ZN (CLOCK_slo__sro_n1471), .A (n_15));
NAND2_X1 CLOCK_slo__sro_c1029 (.ZN (CLOCK_slo__sro_n1470), .A1 (p_1[15]), .A2 (p_0[15]));
OAI21_X4 CLOCK_slo__sro_c1031 (.ZN (CLOCK_slo__sro_n1468), .A (CLOCK_slo__sro_n1470)
    , .B1 (CLOCK_slo__sro_n1471), .B2 (CLOCK_slo__mro_n1886));
XNOR2_X1 CLOCK_slo__sro_c1032 (.ZN (CLOCK_slo__sro_n1467), .A (p_1[15]), .B (p_0[15]));
XNOR2_X1 CLOCK_slo__sro_c1033 (.ZN (p_2[15]), .A (CLOCK_slo__sro_n1467), .B (n_15));
NAND2_X1 CLOCK_slo__sro_c1113 (.ZN (CLOCK_slo__sro_n1550), .A1 (p_1[6]), .A2 (p_0[6]));
NOR2_X1 CLOCK_slo__sro_c1114 (.ZN (CLOCK_slo__sro_n1549), .A1 (p_1[6]), .A2 (p_0[6]));
OAI21_X1 CLOCK_slo__sro_c1115 (.ZN (n_7), .A (CLOCK_slo__sro_n1550), .B1 (CLOCK_slo__sro_n1549), .B2 (CLOCK_slo__sro_n1551));
XNOR2_X1 CLOCK_slo__sro_c1116 (.ZN (CLOCK_slo__sro_n1548), .A (p_1[6]), .B (p_0[6]));
XNOR2_X1 CLOCK_slo__sro_c1117 (.ZN (p_2[6]), .A (CLOCK_slo__sro_n1548), .B (n_6));
NAND2_X1 CLOCK_slo__sro_c1202 (.ZN (CLOCK_slo__sro_n1635), .A1 (n_9), .A2 (p_0[9]));
AOI22_X1 CLOCK_slo__sro_c1203 (.ZN (CLOCK_slo__sro_n1634), .A1 (n_9), .A2 (p_1[9])
    , .B1 (p_1[9]), .B2 (p_0[9]));
NAND2_X1 CLOCK_slo__sro_c1204 (.ZN (n_10), .A1 (CLOCK_slo__sro_n1634), .A2 (CLOCK_slo__sro_n1635));
XNOR2_X1 CLOCK_slo__sro_c1205 (.ZN (CLOCK_slo__sro_n1633), .A (p_1[9]), .B (p_0[9]));
XNOR2_X1 CLOCK_slo__sro_c1206 (.ZN (p_2[9]), .A (CLOCK_slo__sro_n1633), .B (n_9));
NAND2_X1 CLOCK_slo__sro_c1156 (.ZN (CLOCK_slo__sro_n1594), .A1 (p_1[10]), .A2 (p_0[10]));
OAI21_X1 CLOCK_slo__sro_c1157 (.ZN (CLOCK_slo__sro_n1593), .A (n_10), .B1 (p_1[10]), .B2 (p_0[10]));
NAND2_X1 CLOCK_slo__sro_c1158 (.ZN (n_11), .A1 (CLOCK_slo__sro_n1593), .A2 (CLOCK_slo__sro_n1594));
XNOR2_X1 CLOCK_slo__sro_c1159 (.ZN (CLOCK_slo__sro_n1592), .A (p_1[10]), .B (p_0[10]));
XNOR2_X1 CLOCK_slo__sro_c1160 (.ZN (p_2[10]), .A (CLOCK_slo__sro_n1592), .B (n_10));
OAI21_X1 CLOCK_slo__sro_c1350 (.ZN (n_18), .A (CLOCK_slo__sro_n1807), .B1 (CLOCK_slo__sro_n1806), .B2 (CLOCK_slo__sro_n1808));
OAI21_X1 CLOCK_slo__sro_c1330 (.ZN (n_30), .A (slo__sro_n600), .B1 (slo__sro_n601), .B2 (slo__sro_n599));
NOR2_X1 CLOCK_slo__sro_c1349 (.ZN (CLOCK_slo__sro_n1806), .A1 (p_1[17]), .A2 (p_0[17]));
XNOR2_X1 CLOCK_slo__sro_c1351 (.ZN (CLOCK_slo__sro_n1805), .A (p_1[17]), .B (p_0[17]));
XNOR2_X1 CLOCK_slo__sro_c1352 (.ZN (p_2[17]), .A (CLOCK_slo__sro_n1805), .B (n_17));

endmodule //datapath__0_212

module datapath__0_211 (drc_ipoPP_0, Multiplier, p_0, p_1);

output [31:0] p_1;
input [31:0] Multiplier;
input [31:0] p_0;
input drc_ipoPP_0;
wire slo__sro_n529;
wire CLOCK_slo__sro_n1623;
wire n_1;
wire n_2;
wire n_3;
wire n_4;
wire n_5;
wire n_6;
wire n_7;
wire n_8;
wire n_9;
wire n_11;
wire n_12;
wire n_13;
wire n_14;
wire n_15;
wire CLOCK_slo__sro_n1619;
wire CLOCK_slo__mro_n1736;
wire n_20;
wire n_21;
wire n_22;
wire n_23;
wire n_27;
wire n_30;
wire n_32;
wire n_0;
wire n_34;
wire n_33;
wire n_31;
wire slo__sro_n819;
wire slo__sro_n818;
wire slo__sro_n61;
wire slo__sro_n62;
wire slo__sro_n63;
wire slo__sro_n64;
wire slo__sro_n89;
wire slo__sro_n90;
wire slo__sro_n91;
wire slo__sro_n92;
wire slo__sro_n93;
wire slo__sro_n106;
wire slo__sro_n107;
wire slo__sro_n108;
wire slo__sro_n109;
wire slo__sro_n123;
wire slo__sro_n124;
wire slo__sro_n125;
wire slo__sro_n126;
wire slo__sro_n151;
wire slo__sro_n152;
wire slo__sro_n153;
wire slo__sro_n235;
wire slo__sro_n236;
wire slo__sro_n237;
wire slo__sro_n247;
wire slo__sro_n248;
wire slo__sro_n249;
wire slo__sro_n250;
wire slo__sro_n262;
wire slo__sro_n263;
wire slo__sro_n264;
wire slo__sro_n265;
wire slo__sro_n266;
wire slo__sro_n282;
wire slo__sro_n284;
wire slo__sro_n301;
wire slo__sro_n302;
wire slo__sro_n303;
wire slo__sro_n304;
wire slo__sro_n420;
wire CLOCK_slo__sro_n1813;
wire slo__sro_n421;
wire slo__sro_n422;
wire slo__sro_n423;
wire slo__sro_n447;
wire slo__sro_n448;
wire slo__sro_n449;
wire slo__sro_n450;
wire slo__sro_n451;
wire slo__sro_n530;
wire slo__sro_n531;
wire slo__sro_n532;
wire slo__sro_n542;
wire slo__sro_n543;
wire slo__sro_n544;
wire slo__sro_n545;
wire slo__sro_n835;
wire slo__sro_n820;
wire slo__mro_n777;
wire CLOCK_slo__sro_n1749;
wire slo__sro_n834;
wire slo__sro_n821;
wire slo__sro_n836;
wire slo__sro_n837;
wire CLOCK_slo__sro_n1691;
wire CLOCK_slo__sro_n1689;
wire CLOCK_slo__sro_n1690;
wire slo__sro_n889;
wire slo__sro_n890;
wire slo__sro_n891;
wire slo__sro_n892;
wire slo__sro_n893;
wire CLOCK_slo__sro_n1620;
wire CLOCK_slo__sro_n1621;
wire CLOCK_slo__sro_n1622;
wire slo__sro_n1201;
wire slo__sro_n1202;
wire slo__sro_n1203;
wire slo__sro_n1204;
wire CLOCK_slo__sro_n1692;
wire CLOCK_slo__mro_n1704;
wire CLOCK_slo__sro_n1750;
wire CLOCK_slo__sro_n1751;
wire CLOCK_slo__sro_n1752;
wire CLOCK_slo__sro_n1775;
wire CLOCK_slo__sro_n1776;
wire CLOCK_slo__sro_n1777;
wire CLOCK_slo__mro_n1788;
wire CLOCK_slo__mro_n1789;
wire CLOCK_slo__mro_n1790;
wire CLOCK_slo__mro_n1791;
wire CLOCK_slo__sro_n1825;
wire CLOCK_slo__sro_n1826;
wire CLOCK_slo__sro_n1827;
wire CLOCK_slo__sro_n1828;
wire CLOCK_slo__xsl_n2029;


INV_X1 i_36 (.ZN (n_34), .A (Multiplier[30]));
INV_X2 i_35 (.ZN (n_33), .A (p_0[30]));
INV_X1 i_34 (.ZN (n_32), .A (n_30));
OAI33_X1 i_33 (.ZN (n_31), .A1 (n_32), .A2 (p_0[30]), .A3 (n_34), .B1 (n_30), .B2 (n_33), .B3 (Multiplier[30]));
XOR2_X1 i_32 (.Z (p_1[31]), .A (Multiplier[31]), .B (n_31));
OAI22_X1 i_31 (.ZN (n_0), .A1 (n_34), .A2 (p_0[30]), .B1 (n_33), .B2 (Multiplier[30]));
XNOR2_X1 i_0 (.ZN (p_1[30]), .A (n_0), .B (n_32));
INV_X1 slo__sro_c332 (.ZN (slo__sro_n451), .A (slo__sro_n834));
NAND2_X1 slo__sro_c390 (.ZN (slo__sro_n531), .A1 (p_0[3]), .A2 (Multiplier[3]));
OAI21_X1 CLOCK_slo__sro_c1195 (.ZN (n_6), .A (CLOCK_slo__sro_n1691), .B1 (CLOCK_slo__sro_n1690), .B2 (CLOCK_slo__sro_n1692));
FA_X1 i_27 (.CO (n_27), .S (p_1[26]), .A (Multiplier[26]), .B (p_0[26]), .CI (slo__sro_n107));
INV_X1 slo__sro_c59 (.ZN (slo__sro_n126), .A (n_7));
INV_X1 slo__sro_c231 (.ZN (slo__sro_n304), .A (n_21));
INV_X2 slo__sro_c31 (.ZN (slo__sro_n93), .A (CLOCK_slo__sro_n1620));
INV_X1 slo__sro_c389 (.ZN (slo__sro_n532), .A (n_3));
FA_X1 i_21 (.CO (n_21), .S (p_1[20]), .A (Multiplier[20]), .B (p_0[20]), .CI (n_20));
INV_X1 slo__sro_c165 (.ZN (slo__sro_n237), .A (p_0[8]));
INV_X1 CLOCK_slo__sro_c1192 (.ZN (CLOCK_slo__sro_n1692), .A (n_5));
NAND2_X1 slo__sro_c211 (.ZN (slo__sro_n284), .A1 (p_0[24]), .A2 (Multiplier[24]));
NAND3_X2 CLOCK_slo__sro_c1117 (.ZN (CLOCK_slo__sro_n1620), .A1 (CLOCK_slo__sro_n1621)
    , .A2 (CLOCK_slo__sro_n1622), .A3 (CLOCK_slo__sro_n1623));
INV_X1 slo__sro_c195 (.ZN (slo__sro_n266), .A (slo__sro_n890));
NAND2_X1 CLOCK_slo__sro_c1193 (.ZN (CLOCK_slo__sro_n1691), .A1 (p_0[5]), .A2 (Multiplier[5]));
FA_X1 i_13 (.CO (n_13), .S (p_1[12]), .A (Multiplier[12]), .B (p_0[12]), .CI (n_12));
FA_X1 i_12 (.CO (n_12), .S (p_1[11]), .A (Multiplier[11]), .B (p_0[11]), .CI (n_11));
INV_X1 CLOCK_slo__mro_c1295 (.ZN (CLOCK_slo__mro_n1791), .A (Multiplier[8]));
INV_X1 slo__sro_c179 (.ZN (slo__sro_n250), .A (n_14));
NAND2_X1 slo__sro_c86 (.ZN (slo__sro_n153), .A1 (slo__sro_n90), .A2 (Multiplier[19]));
INV_X1 slo__sro_c633 (.ZN (slo__sro_n837), .A (n_27));
XNOR2_X2 CLOCK_slo__mro_c1214 (.ZN (CLOCK_slo__mro_n1704), .A (slo__sro_n61), .B (Multiplier[24]));
FA_X1 i_5 (.CO (n_5), .S (p_1[4]), .A (Multiplier[4]), .B (p_0[4]), .CI (n_4));
INV_X1 slo__sro_c403 (.ZN (slo__sro_n545), .A (p_0[1]));
FA_X1 i_3 (.CO (n_3), .S (p_1[2]), .A (Multiplier[2]), .B (p_0[2]), .CI (n_2));
INV_X1 slo__sro_c617 (.ZN (slo__sro_n821), .A (p_0[6]));
HA_X1 i_1 (.CO (n_1), .S (p_1[0]), .A (Multiplier[0]), .B (p_0[0]));
INV_X2 slo__sro_c4 (.ZN (slo__sro_n64), .A (n_23));
NAND2_X1 slo__sro_c5 (.ZN (slo__sro_n63), .A1 (p_0[23]), .A2 (Multiplier[23]));
NOR2_X2 slo__sro_c6 (.ZN (slo__sro_n62), .A1 (p_0[23]), .A2 (Multiplier[23]));
OAI21_X2 slo__sro_c7 (.ZN (slo__sro_n61), .A (slo__sro_n63), .B1 (slo__sro_n62), .B2 (slo__sro_n64));
NOR2_X1 slo__sro_c619 (.ZN (slo__sro_n819), .A1 (n_6), .A2 (Multiplier[6]));
OAI21_X2 slo__sro_c620 (.ZN (n_7), .A (slo__sro_n820), .B1 (slo__sro_n821), .B2 (slo__sro_n819));
NAND2_X1 slo__sro_c32 (.ZN (slo__sro_n92), .A1 (p_0[18]), .A2 (Multiplier[18]));
NOR2_X2 slo__sro_c33 (.ZN (slo__sro_n91), .A1 (p_0[18]), .A2 (Multiplier[18]));
OAI21_X2 slo__sro_c34 (.ZN (slo__sro_n90), .A (slo__sro_n92), .B1 (slo__sro_n93), .B2 (slo__sro_n91));
XNOR2_X1 slo__sro_c35 (.ZN (slo__sro_n89), .A (p_0[18]), .B (Multiplier[18]));
XNOR2_X1 slo__sro_c36 (.ZN (p_1[18]), .A (slo__sro_n89), .B (CLOCK_slo__sro_n1620));
NAND2_X1 slo__sro_c46 (.ZN (slo__sro_n109), .A1 (p_0[25]), .A2 (Multiplier[25]));
NOR2_X1 slo__sro_c47 (.ZN (slo__sro_n108), .A1 (p_0[25]), .A2 (Multiplier[25]));
OAI21_X2 slo__sro_c48 (.ZN (slo__sro_n107), .A (slo__sro_n109), .B1 (slo__sro_n108), .B2 (slo__sro_n282));
XNOR2_X2 slo__sro_c49 (.ZN (slo__sro_n106), .A (p_0[25]), .B (Multiplier[25]));
XNOR2_X2 slo__sro_c50 (.ZN (p_1[25]), .A (slo__sro_n106), .B (CLOCK_slo__xsl_n2029));
NAND2_X1 slo__sro_c60 (.ZN (slo__sro_n125), .A1 (p_0[7]), .A2 (Multiplier[7]));
NOR2_X2 slo__sro_c61 (.ZN (slo__sro_n124), .A1 (p_0[7]), .A2 (drc_ipoPP_0));
OAI21_X2 slo__sro_c62 (.ZN (n_8), .A (slo__sro_n125), .B1 (slo__sro_n126), .B2 (slo__sro_n124));
XNOR2_X2 slo__sro_c63 (.ZN (slo__sro_n123), .A (p_0[7]), .B (Multiplier[7]));
XNOR2_X2 slo__sro_c64 (.ZN (p_1[7]), .A (slo__sro_n123), .B (n_7));
OAI21_X1 slo__sro_c87 (.ZN (slo__sro_n152), .A (p_0[19]), .B1 (slo__sro_n90), .B2 (Multiplier[19]));
NAND2_X1 slo__sro_c88 (.ZN (n_20), .A1 (slo__sro_n152), .A2 (slo__sro_n153));
XNOR2_X2 slo__sro_c89 (.ZN (slo__sro_n151), .A (slo__sro_n90), .B (Multiplier[19]));
XNOR2_X2 slo__sro_c90 (.ZN (p_1[19]), .A (slo__sro_n151), .B (p_0[19]));
NAND2_X1 slo__sro_c166 (.ZN (slo__sro_n236), .A1 (n_8), .A2 (Multiplier[8]));
NOR2_X2 slo__sro_c167 (.ZN (slo__sro_n235), .A1 (n_8), .A2 (Multiplier[8]));
OAI21_X2 slo__sro_c168 (.ZN (n_9), .A (slo__sro_n236), .B1 (slo__sro_n237), .B2 (slo__sro_n235));
OAI21_X1 CLOCK_slo__sro_c1319 (.ZN (CLOCK_slo__sro_n1813), .A (slo__sro_n61), .B1 (p_0[24]), .B2 (Multiplier[24]));
NAND2_X1 CLOCK_slo__sro_c1329 (.ZN (CLOCK_slo__sro_n1828), .A1 (p_0[22]), .A2 (Multiplier[22]));
NAND2_X1 slo__sro_c180 (.ZN (slo__sro_n249), .A1 (p_0[14]), .A2 (Multiplier[14]));
NOR2_X1 slo__sro_c181 (.ZN (slo__sro_n248), .A1 (p_0[14]), .A2 (Multiplier[14]));
OAI21_X2 slo__sro_c182 (.ZN (n_15), .A (slo__sro_n249), .B1 (slo__sro_n250), .B2 (slo__sro_n248));
XNOR2_X1 slo__sro_c183 (.ZN (slo__sro_n247), .A (p_0[14]), .B (Multiplier[14]));
XNOR2_X1 slo__sro_c184 (.ZN (p_1[14]), .A (slo__sro_n247), .B (n_14));
NAND2_X1 slo__sro_c196 (.ZN (slo__sro_n265), .A1 (p_0[16]), .A2 (Multiplier[16]));
NOR2_X2 slo__sro_c197 (.ZN (slo__sro_n264), .A1 (p_0[16]), .A2 (Multiplier[16]));
OAI21_X2 slo__sro_c198 (.ZN (slo__sro_n263), .A (slo__sro_n265), .B1 (slo__sro_n264), .B2 (slo__sro_n266));
XNOR2_X2 slo__sro_c199 (.ZN (slo__sro_n262), .A (p_0[16]), .B (Multiplier[16]));
XNOR2_X1 slo__sro_c200 (.ZN (p_1[16]), .A (slo__sro_n262), .B (slo__sro_n890));
INV_X1 CLOCK_slo__xsl_c1511 (.ZN (CLOCK_slo__xsl_n2029), .A (slo__sro_n282));
XNOR2_X2 CLOCK_slo__mro_c1247 (.ZN (CLOCK_slo__mro_n1736), .A (p_0[27]), .B (Multiplier[27]));
XNOR2_X2 CLOCK_slo__mro_c1248 (.ZN (p_1[27]), .A (CLOCK_slo__mro_n1736), .B (n_27));
NAND2_X1 slo__sro_c232 (.ZN (slo__sro_n303), .A1 (p_0[21]), .A2 (Multiplier[21]));
NOR2_X2 slo__sro_c233 (.ZN (slo__sro_n302), .A1 (p_0[21]), .A2 (Multiplier[21]));
OAI21_X2 slo__sro_c234 (.ZN (n_22), .A (slo__sro_n303), .B1 (slo__sro_n304), .B2 (slo__sro_n302));
XNOR2_X2 slo__sro_c235 (.ZN (slo__sro_n301), .A (p_0[21]), .B (Multiplier[21]));
XNOR2_X1 slo__sro_c236 (.ZN (p_1[21]), .A (slo__sro_n301), .B (n_21));
INV_X1 slo__sro_c303 (.ZN (slo__sro_n423), .A (slo__sro_n448));
NAND2_X1 slo__sro_c304 (.ZN (slo__sro_n422), .A1 (p_0[29]), .A2 (Multiplier[29]));
NOR2_X1 slo__sro_c305 (.ZN (slo__sro_n421), .A1 (p_0[29]), .A2 (Multiplier[29]));
OAI21_X1 slo__sro_c306 (.ZN (n_30), .A (slo__sro_n422), .B1 (slo__sro_n423), .B2 (slo__sro_n421));
XNOR2_X1 slo__sro_c307 (.ZN (slo__sro_n420), .A (p_0[29]), .B (Multiplier[29]));
XNOR2_X1 slo__sro_c308 (.ZN (p_1[29]), .A (slo__sro_n420), .B (slo__sro_n448));
NAND2_X1 slo__sro_c333 (.ZN (slo__sro_n450), .A1 (p_0[28]), .A2 (Multiplier[28]));
NOR2_X1 slo__sro_c334 (.ZN (slo__sro_n449), .A1 (p_0[28]), .A2 (Multiplier[28]));
OAI21_X2 slo__sro_c335 (.ZN (slo__sro_n448), .A (slo__sro_n450), .B1 (slo__sro_n449), .B2 (slo__sro_n451));
XNOR2_X2 slo__sro_c336 (.ZN (slo__sro_n447), .A (p_0[28]), .B (Multiplier[28]));
XNOR2_X1 slo__sro_c337 (.ZN (p_1[28]), .A (slo__sro_n447), .B (slo__sro_n834));
NOR2_X1 slo__sro_c391 (.ZN (slo__sro_n530), .A1 (p_0[3]), .A2 (Multiplier[3]));
OAI21_X1 slo__sro_c392 (.ZN (n_4), .A (slo__sro_n531), .B1 (slo__sro_n532), .B2 (slo__sro_n530));
XNOR2_X1 slo__sro_c393 (.ZN (slo__sro_n529), .A (p_0[3]), .B (Multiplier[3]));
XNOR2_X1 slo__sro_c394 (.ZN (p_1[3]), .A (slo__sro_n529), .B (n_3));
NAND2_X1 slo__sro_c404 (.ZN (slo__sro_n544), .A1 (n_1), .A2 (Multiplier[1]));
NOR2_X1 slo__sro_c405 (.ZN (slo__sro_n543), .A1 (n_1), .A2 (Multiplier[1]));
OAI21_X1 slo__sro_c406 (.ZN (n_2), .A (slo__sro_n544), .B1 (slo__sro_n545), .B2 (slo__sro_n543));
XNOR2_X1 slo__sro_c407 (.ZN (slo__sro_n542), .A (n_1), .B (Multiplier[1]));
XNOR2_X1 slo__sro_c408 (.ZN (p_1[1]), .A (slo__sro_n542), .B (p_0[1]));
NAND2_X1 slo__sro_c618 (.ZN (slo__sro_n820), .A1 (n_6), .A2 (Multiplier[6]));
XNOR2_X1 slo__sro_c621 (.ZN (slo__sro_n818), .A (n_6), .B (Multiplier[6]));
XNOR2_X2 slo__mro_c578 (.ZN (slo__mro_n777), .A (p_0[23]), .B (Multiplier[23]));
XNOR2_X2 slo__mro_c579 (.ZN (p_1[23]), .A (slo__mro_n777), .B (n_23));
NAND2_X1 slo__sro_c634 (.ZN (slo__sro_n836), .A1 (p_0[27]), .A2 (Multiplier[27]));
NOR2_X1 slo__sro_c635 (.ZN (slo__sro_n835), .A1 (p_0[27]), .A2 (Multiplier[27]));
OAI21_X1 slo__sro_c636 (.ZN (slo__sro_n834), .A (slo__sro_n836), .B1 (slo__sro_n837), .B2 (slo__sro_n835));
NAND2_X1 CLOCK_slo__sro_c1260 (.ZN (CLOCK_slo__sro_n1752), .A1 (n_9), .A2 (Multiplier[9]));
XNOR2_X1 slo__sro_c622 (.ZN (p_1[6]), .A (slo__sro_n818), .B (p_0[6]));
OAI21_X1 CLOCK_slo__sro_c1261 (.ZN (CLOCK_slo__sro_n1751), .A (p_0[9]), .B1 (n_9), .B2 (Multiplier[9]));
XNOR2_X1 CLOCK_slo__sro_c1196 (.ZN (CLOCK_slo__sro_n1689), .A (p_0[5]), .B (Multiplier[5]));
NOR2_X1 CLOCK_slo__sro_c1194 (.ZN (CLOCK_slo__sro_n1690), .A1 (p_0[5]), .A2 (Multiplier[5]));
NAND2_X1 CLOCK_slo__sro_c1114 (.ZN (CLOCK_slo__sro_n1623), .A1 (p_0[17]), .A2 (Multiplier[17]));
NAND2_X1 CLOCK_slo__sro_c1115 (.ZN (CLOCK_slo__sro_n1622), .A1 (slo__sro_n263), .A2 (Multiplier[17]));
NAND2_X1 CLOCK_slo__sro_c1116 (.ZN (CLOCK_slo__sro_n1621), .A1 (slo__sro_n263), .A2 (p_0[17]));
INV_X1 slo__sro_c679 (.ZN (slo__sro_n893), .A (n_15));
NAND2_X1 slo__sro_c680 (.ZN (slo__sro_n892), .A1 (p_0[15]), .A2 (Multiplier[15]));
NOR2_X1 slo__sro_c681 (.ZN (slo__sro_n891), .A1 (p_0[15]), .A2 (Multiplier[15]));
OAI21_X1 slo__sro_c682 (.ZN (slo__sro_n890), .A (slo__sro_n892), .B1 (slo__sro_n891), .B2 (slo__sro_n893));
XNOR2_X1 slo__sro_c683 (.ZN (slo__sro_n889), .A (p_0[15]), .B (Multiplier[15]));
XNOR2_X1 slo__sro_c684 (.ZN (p_1[15]), .A (slo__sro_n889), .B (n_15));
XNOR2_X1 CLOCK_slo__sro_c1118 (.ZN (CLOCK_slo__sro_n1619), .A (p_0[17]), .B (Multiplier[17]));
XNOR2_X1 CLOCK_slo__sro_c1119 (.ZN (p_1[17]), .A (CLOCK_slo__sro_n1619), .B (slo__sro_n263));
INV_X1 slo__sro_c851 (.ZN (slo__sro_n1204), .A (n_13));
NAND2_X1 slo__sro_c852 (.ZN (slo__sro_n1203), .A1 (p_0[13]), .A2 (Multiplier[13]));
NOR2_X1 slo__sro_c853 (.ZN (slo__sro_n1202), .A1 (p_0[13]), .A2 (Multiplier[13]));
OAI21_X2 slo__sro_c854 (.ZN (n_14), .A (slo__sro_n1203), .B1 (slo__sro_n1204), .B2 (slo__sro_n1202));
XNOR2_X1 slo__sro_c855 (.ZN (slo__sro_n1201), .A (p_0[13]), .B (Multiplier[13]));
XNOR2_X1 slo__sro_c856 (.ZN (p_1[13]), .A (slo__sro_n1201), .B (n_13));
XNOR2_X1 CLOCK_slo__sro_c1197 (.ZN (p_1[5]), .A (CLOCK_slo__sro_n1689), .B (n_5));
XNOR2_X2 CLOCK_slo__mro_c1215 (.ZN (p_1[24]), .A (p_0[24]), .B (CLOCK_slo__mro_n1704));
NAND2_X1 CLOCK_slo__sro_c1262 (.ZN (CLOCK_slo__sro_n1750), .A1 (CLOCK_slo__sro_n1752), .A2 (CLOCK_slo__sro_n1751));
XNOR2_X1 CLOCK_slo__sro_c1263 (.ZN (CLOCK_slo__sro_n1749), .A (p_0[9]), .B (Multiplier[9]));
XNOR2_X1 CLOCK_slo__sro_c1264 (.ZN (p_1[9]), .A (CLOCK_slo__sro_n1749), .B (n_9));
NAND2_X1 CLOCK_slo__sro_c1283 (.ZN (CLOCK_slo__sro_n1777), .A1 (CLOCK_slo__sro_n1750), .A2 (Multiplier[10]));
AOI22_X1 CLOCK_slo__sro_c1284 (.ZN (CLOCK_slo__sro_n1776), .A1 (CLOCK_slo__sro_n1750)
    , .A2 (p_0[10]), .B1 (p_0[10]), .B2 (Multiplier[10]));
NAND2_X1 CLOCK_slo__sro_c1285 (.ZN (n_11), .A1 (CLOCK_slo__sro_n1776), .A2 (CLOCK_slo__sro_n1777));
XNOR2_X1 CLOCK_slo__sro_c1286 (.ZN (CLOCK_slo__sro_n1775), .A (p_0[10]), .B (Multiplier[10]));
XNOR2_X1 CLOCK_slo__sro_c1287 (.ZN (p_1[10]), .A (CLOCK_slo__sro_n1775), .B (CLOCK_slo__sro_n1750));
OAI21_X1 CLOCK_slo__mro_c1296 (.ZN (CLOCK_slo__mro_n1790), .A (slo__sro_n125), .B1 (slo__sro_n124), .B2 (slo__sro_n126));
INV_X1 CLOCK_slo__mro_c1297 (.ZN (CLOCK_slo__mro_n1789), .A (CLOCK_slo__mro_n1790));
XNOR2_X2 CLOCK_slo__mro_c1298 (.ZN (CLOCK_slo__mro_n1788), .A (p_0[8]), .B (CLOCK_slo__mro_n1791));
XNOR2_X2 CLOCK_slo__mro_c1299 (.ZN (p_1[8]), .A (CLOCK_slo__mro_n1788), .B (CLOCK_slo__mro_n1789));
NAND2_X2 CLOCK_slo__sro_c1330 (.ZN (CLOCK_slo__sro_n1827), .A1 (n_22), .A2 (Multiplier[22]));
NAND2_X1 CLOCK_slo__sro_c1331 (.ZN (CLOCK_slo__sro_n1826), .A1 (n_22), .A2 (p_0[22]));
NAND3_X2 CLOCK_slo__sro_c1332 (.ZN (n_23), .A1 (CLOCK_slo__sro_n1827), .A2 (CLOCK_slo__sro_n1826), .A3 (CLOCK_slo__sro_n1828));
XNOR2_X2 CLOCK_slo__sro_c1333 (.ZN (CLOCK_slo__sro_n1825), .A (p_0[22]), .B (Multiplier[22]));
XNOR2_X1 CLOCK_slo__sro_c1334 (.ZN (p_1[22]), .A (CLOCK_slo__sro_n1825), .B (n_22));
AND2_X1 CLOCK_slo__xsl_c1514 (.ZN (slo__sro_n282), .A1 (CLOCK_slo__sro_n1813), .A2 (slo__sro_n284));

endmodule //datapath__0_211

module datapath__0_207 (p_0, p_1, p_2);

output [31:0] p_2;
input [31:0] p_0;
input [31:0] p_1;
wire CLOCK_slo__sro_n1086;
wire n_1;
wire n_2;
wire n_3;
wire n_4;
wire n_5;
wire n_6;
wire n_7;
wire n_8;
wire n_9;
wire n_10;
wire n_11;
wire n_12;
wire n_13;
wire n_14;
wire n_15;
wire CLOCK_slo__sro_n1441;
wire n_18;
wire n_19;
wire n_20;
wire n_21;
wire n_22;
wire n_23;
wire slo__sro_n470;
wire n_25;
wire n_26;
wire n_27;
wire n_28;
wire n_29;
wire n_30;
wire n_32;
wire n_0;
wire n_34;
wire n_33;
wire slo__sro_n129;
wire slo__sro_n130;
wire slo__sro_n131;
wire slo__sro_n132;
wire slo__sro_n273;
wire slo__sro_n274;
wire slo__sro_n275;
wire slo__sro_n276;
wire slo__sro_n299;
wire slo__sro_n300;
wire slo__sro_n301;
wire slo__sro_n302;
wire slo__sro_n170;
wire slo__sro_n171;
wire slo__sro_n172;
wire slo__sro_n426;
wire slo__sro_n427;
wire slo__sro_n428;
wire slo__sro_n429;
wire slo__sro_n439;
wire slo__sro_n224;
wire slo__sro_n225;
wire slo__sro_n226;
wire slo__sro_n227;
wire slo__sro_n440;
wire slo__sro_n441;
wire slo__sro_n442;
wire slo__sro_n443;
wire slo__sro_n471;
wire slo__sro_n472;
wire slo__sro_n473;
wire slo__sro_n474;
wire slo__sro_n496;
wire slo__sro_n497;
wire slo__sro_n498;
wire slo__sro_n499;
wire CLOCK_slo__sro_n1054;
wire slo__sro_n536;
wire slo__sro_n537;
wire slo__sro_n538;
wire slo__sro_n539;
wire CLOCK_slo__sro_n1087;
wire CLOCK_slo__mro_n1064;
wire CLOCK_slo__sro_n1051;
wire CLOCK_slo__sro_n1052;
wire CLOCK_slo__sro_n1053;
wire slo__sro_n564;
wire slo__sro_n565;
wire slo__sro_n566;
wire slo__sro_n567;
wire CLOCK_slo__sro_n1088;
wire CLOCK_slo__sro_n1089;
wire CLOCK_slo__sro_n1150;
wire CLOCK_slo__sro_n1151;
wire CLOCK_slo__sro_n1152;
wire CLOCK_slo__sro_n1153;
wire CLOCK_slo__sro_n1246;
wire CLOCK_slo__sro_n1247;
wire CLOCK_slo__sro_n1248;
wire CLOCK_slo__sro_n1249;
wire CLOCK_slo__sro_n1250;
wire CLOCK_slo__sro_n1442;
wire CLOCK_slo__sro_n1443;


INV_X1 i_36 (.ZN (n_34), .A (p_0[30]));
INV_X1 i_35 (.ZN (n_33), .A (p_1[30]));
INV_X1 i_34 (.ZN (n_32), .A (n_30));
INV_X1 slo__sro_c378 (.ZN (slo__sro_n499), .A (n_27));
XOR2_X1 i_32 (.Z (p_2[31]), .A (p_0[31]), .B (slo__sro_n470));
OAI22_X1 i_31 (.ZN (n_0), .A1 (n_34), .A2 (p_1[30]), .B1 (p_0[30]), .B2 (n_33));
XNOR2_X1 i_0 (.ZN (p_2[30]), .A (n_32), .B (n_0));
FA_X1 i_30 (.CO (n_30), .S (p_2[29]), .A (p_0[29]), .B (p_1[29]), .CI (n_29));
FA_X1 i_29 (.CO (n_29), .S (p_2[28]), .A (p_0[28]), .B (p_1[28]), .CI (n_28));
XNOR2_X1 CLOCK_slo__sro_c738 (.ZN (p_2[9]), .A (CLOCK_slo__sro_n1051), .B (n_9));
OAI21_X2 CLOCK_slo__sro_c975 (.ZN (n_5), .A (slo__sro_n171), .B1 (slo__sro_n170), .B2 (slo__sro_n172));
XNOR2_X1 CLOCK_slo__sro_c737 (.ZN (CLOCK_slo__sro_n1051), .A (p_1[9]), .B (p_0[9]));
FA_X1 i_25 (.CO (n_25), .S (p_2[24]), .A (p_0[24]), .B (p_1[24]), .CI (slo__sro_n440));
INV_X1 slo__sro_c353 (.ZN (slo__sro_n474), .A (n_30));
FA_X1 i_23 (.CO (n_23), .S (p_2[22]), .A (p_0[22]), .B (p_1[22]), .CI (n_22));
INV_X1 slo__sro_c329 (.ZN (slo__sro_n443), .A (n_23));
FA_X1 i_21 (.CO (n_21), .S (p_2[20]), .A (p_0[20]), .B (p_1[20]), .CI (n_20));
OAI21_X1 slo__sro_c332 (.ZN (slo__sro_n440), .A (slo__sro_n442), .B1 (slo__sro_n443), .B2 (slo__sro_n441));
FA_X1 i_19 (.CO (n_19), .S (p_2[18]), .A (p_0[18]), .B (p_1[18]), .CI (n_18));
INV_X1 slo__sro_c232 (.ZN (slo__sro_n302), .A (n_11));
INV_X1 CLOCK_slo__sro_c840 (.ZN (CLOCK_slo__sro_n1153), .A (p_1[26]));
NAND2_X1 CLOCK_slo__sro_c1124 (.ZN (CLOCK_slo__sro_n1443), .A1 (n_1), .A2 (p_0[1]));
XNOR2_X1 CLOCK_slo__sro_c768 (.ZN (CLOCK_slo__sro_n1086), .A (p_1[16]), .B (p_0[16]));
FA_X1 i_14 (.CO (n_14), .S (p_2[13]), .A (p_0[13]), .B (p_1[13]), .CI (n_13));
FA_X1 i_13 (.CO (n_13), .S (p_2[12]), .A (p_0[12]), .B (p_1[12]), .CI (n_12));
INV_X1 slo__sro_c315 (.ZN (slo__sro_n429), .A (n_21));
INV_X1 slo__sro_c205 (.ZN (slo__sro_n276), .A (CLOCK_slo__sro_n1087));
XNOR2_X2 CLOCK_slo__mro_c747 (.ZN (CLOCK_slo__mro_n1064), .A (p_1[4]), .B (p_0[4]));
FA_X1 i_9 (.CO (n_9), .S (p_2[8]), .A (p_0[8]), .B (p_1[8]), .CI (n_8));
FA_X1 i_8 (.CO (n_8), .S (p_2[7]), .A (p_0[7]), .B (p_1[7]), .CI (n_7));
FA_X1 i_7 (.CO (n_7), .S (p_2[6]), .A (p_0[6]), .B (p_1[6]), .CI (n_6));
FA_X1 i_6 (.CO (n_6), .S (p_2[5]), .A (p_0[5]), .B (p_1[5]), .CI (n_5));
NOR2_X1 slo__sro_c317 (.ZN (slo__sro_n427), .A1 (p_1[21]), .A2 (p_0[21]));
FA_X1 i_4 (.CO (n_4), .S (p_2[3]), .A (p_0[3]), .B (p_1[3]), .CI (n_3));
FA_X1 i_3 (.CO (n_3), .S (p_2[2]), .A (p_0[2]), .B (p_1[2]), .CI (n_2));
HA_X1 i_1 (.CO (n_1), .S (p_2[0]), .A (p_0[0]), .B (p_1[0]));
INV_X1 slo__sro_c66 (.ZN (slo__sro_n132), .A (n_10));
NAND2_X1 slo__sro_c67 (.ZN (slo__sro_n131), .A1 (p_1[10]), .A2 (p_0[10]));
NOR2_X1 slo__sro_c68 (.ZN (slo__sro_n130), .A1 (p_1[10]), .A2 (p_0[10]));
OAI21_X2 slo__sro_c69 (.ZN (n_11), .A (slo__sro_n131), .B1 (slo__sro_n132), .B2 (slo__sro_n130));
XNOR2_X1 slo__sro_c70 (.ZN (slo__sro_n129), .A (p_1[10]), .B (p_0[10]));
XNOR2_X1 slo__sro_c71 (.ZN (p_2[10]), .A (n_10), .B (slo__sro_n129));
NAND2_X1 slo__sro_c206 (.ZN (slo__sro_n275), .A1 (p_1[17]), .A2 (p_0[17]));
NOR2_X1 slo__sro_c207 (.ZN (slo__sro_n274), .A1 (p_1[17]), .A2 (p_0[17]));
OAI21_X1 slo__sro_c208 (.ZN (n_18), .A (slo__sro_n275), .B1 (slo__sro_n276), .B2 (slo__sro_n274));
XNOR2_X1 slo__sro_c209 (.ZN (slo__sro_n273), .A (p_1[17]), .B (p_0[17]));
XNOR2_X1 slo__sro_c210 (.ZN (p_2[17]), .A (slo__sro_n273), .B (CLOCK_slo__sro_n1087));
NAND2_X1 slo__sro_c233 (.ZN (slo__sro_n301), .A1 (p_1[11]), .A2 (p_0[11]));
NOR2_X1 slo__sro_c234 (.ZN (slo__sro_n300), .A1 (p_1[11]), .A2 (p_0[11]));
OAI21_X1 slo__sro_c235 (.ZN (n_12), .A (slo__sro_n301), .B1 (slo__sro_n302), .B2 (slo__sro_n300));
XNOR2_X1 slo__sro_c236 (.ZN (slo__sro_n299), .A (p_1[11]), .B (p_0[11]));
XNOR2_X1 slo__sro_c237 (.ZN (p_2[11]), .A (slo__sro_n299), .B (n_11));
NAND2_X1 slo__sro_c316 (.ZN (slo__sro_n428), .A1 (p_1[21]), .A2 (p_0[21]));
INV_X1 slo__sro_c106 (.ZN (slo__sro_n172), .A (p_1[4]));
NAND2_X1 slo__sro_c107 (.ZN (slo__sro_n171), .A1 (n_4), .A2 (p_0[4]));
NOR2_X2 slo__sro_c108 (.ZN (slo__sro_n170), .A1 (n_4), .A2 (p_0[4]));
NAND2_X1 CLOCK_slo__sro_c765 (.ZN (CLOCK_slo__sro_n1089), .A1 (p_0[16]), .A2 (p_1[16]));
XNOR2_X1 CLOCK_slo__mro_c748 (.ZN (p_2[4]), .A (n_4), .B (CLOCK_slo__mro_n1064));
OAI21_X1 slo__sro_c318 (.ZN (n_22), .A (slo__sro_n428), .B1 (slo__sro_n429), .B2 (slo__sro_n427));
XNOR2_X1 slo__sro_c319 (.ZN (slo__sro_n426), .A (p_1[21]), .B (p_0[21]));
XNOR2_X1 slo__sro_c320 (.ZN (p_2[21]), .A (slo__sro_n426), .B (n_21));
NAND2_X1 slo__sro_c330 (.ZN (slo__sro_n442), .A1 (p_1[23]), .A2 (p_0[23]));
NOR2_X1 slo__sro_c331 (.ZN (slo__sro_n441), .A1 (p_1[23]), .A2 (p_0[23]));
INV_X1 slo__sro_c159 (.ZN (slo__sro_n227), .A (n_19));
NAND2_X1 slo__sro_c160 (.ZN (slo__sro_n226), .A1 (p_1[19]), .A2 (p_0[19]));
NOR2_X1 slo__sro_c161 (.ZN (slo__sro_n225), .A1 (p_1[19]), .A2 (p_0[19]));
OAI21_X1 slo__sro_c162 (.ZN (n_20), .A (slo__sro_n226), .B1 (slo__sro_n227), .B2 (slo__sro_n225));
XNOR2_X1 slo__sro_c163 (.ZN (slo__sro_n224), .A (p_1[19]), .B (p_0[19]));
XNOR2_X1 slo__sro_c164 (.ZN (p_2[19]), .A (slo__sro_n224), .B (n_19));
XNOR2_X1 slo__sro_c333 (.ZN (slo__sro_n439), .A (p_1[23]), .B (p_0[23]));
XNOR2_X1 slo__sro_c334 (.ZN (p_2[23]), .A (slo__sro_n439), .B (n_23));
NOR2_X1 slo__sro_c354 (.ZN (slo__sro_n473), .A1 (n_33), .A2 (p_0[30]));
NAND2_X1 slo__sro_c355 (.ZN (slo__sro_n472), .A1 (slo__sro_n474), .A2 (slo__sro_n473));
OR2_X1 slo__sro_c356 (.ZN (slo__sro_n471), .A1 (p_1[30]), .A2 (n_34));
OAI21_X1 slo__sro_c357 (.ZN (slo__sro_n470), .A (slo__sro_n472), .B1 (n_32), .B2 (slo__sro_n471));
NAND2_X1 slo__sro_c379 (.ZN (slo__sro_n498), .A1 (p_1[27]), .A2 (p_0[27]));
NOR2_X1 slo__sro_c380 (.ZN (slo__sro_n497), .A1 (p_1[27]), .A2 (p_0[27]));
OAI21_X1 slo__sro_c381 (.ZN (n_28), .A (slo__sro_n498), .B1 (slo__sro_n497), .B2 (slo__sro_n499));
XNOR2_X1 slo__sro_c382 (.ZN (slo__sro_n496), .A (p_1[27]), .B (p_0[27]));
XNOR2_X1 slo__sro_c383 (.ZN (p_2[27]), .A (slo__sro_n496), .B (n_27));
OAI21_X1 CLOCK_slo__sro_c766 (.ZN (CLOCK_slo__sro_n1088), .A (CLOCK_slo__sro_n1247)
    , .B1 (p_1[16]), .B2 (p_0[16]));
INV_X1 slo__sro_c418 (.ZN (slo__sro_n539), .A (n_14));
NAND2_X1 slo__sro_c419 (.ZN (slo__sro_n538), .A1 (p_1[14]), .A2 (p_0[14]));
NOR2_X1 slo__sro_c420 (.ZN (slo__sro_n537), .A1 (p_1[14]), .A2 (p_0[14]));
OAI21_X2 slo__sro_c421 (.ZN (n_15), .A (slo__sro_n538), .B1 (slo__sro_n539), .B2 (slo__sro_n537));
XNOR2_X1 slo__sro_c422 (.ZN (slo__sro_n536), .A (p_1[14]), .B (p_0[14]));
XNOR2_X1 slo__sro_c423 (.ZN (p_2[14]), .A (slo__sro_n536), .B (n_14));
NAND2_X1 CLOCK_slo__sro_c767 (.ZN (CLOCK_slo__sro_n1087), .A1 (CLOCK_slo__sro_n1088), .A2 (CLOCK_slo__sro_n1089));
INV_X2 CLOCK_slo__sro_c733 (.ZN (CLOCK_slo__sro_n1054), .A (n_9));
NAND2_X1 CLOCK_slo__sro_c734 (.ZN (CLOCK_slo__sro_n1053), .A1 (p_1[9]), .A2 (p_0[9]));
NOR2_X1 CLOCK_slo__sro_c735 (.ZN (CLOCK_slo__sro_n1052), .A1 (p_1[9]), .A2 (p_0[9]));
OAI21_X2 CLOCK_slo__sro_c736 (.ZN (n_10), .A (CLOCK_slo__sro_n1053), .B1 (CLOCK_slo__sro_n1054), .B2 (CLOCK_slo__sro_n1052));
INV_X1 slo__sro_c445 (.ZN (slo__sro_n567), .A (n_25));
NAND2_X1 slo__sro_c446 (.ZN (slo__sro_n566), .A1 (p_1[25]), .A2 (p_0[25]));
NOR2_X1 slo__sro_c447 (.ZN (slo__sro_n565), .A1 (p_1[25]), .A2 (p_0[25]));
OAI21_X2 slo__sro_c448 (.ZN (n_26), .A (slo__sro_n566), .B1 (slo__sro_n567), .B2 (slo__sro_n565));
XNOR2_X1 slo__sro_c449 (.ZN (slo__sro_n564), .A (p_1[25]), .B (p_0[25]));
XNOR2_X1 slo__sro_c450 (.ZN (p_2[25]), .A (slo__sro_n564), .B (n_25));
XNOR2_X1 CLOCK_slo__sro_c769 (.ZN (p_2[16]), .A (CLOCK_slo__sro_n1086), .B (CLOCK_slo__sro_n1247));
NAND2_X1 CLOCK_slo__sro_c841 (.ZN (CLOCK_slo__sro_n1152), .A1 (n_26), .A2 (p_0[26]));
NOR2_X1 CLOCK_slo__sro_c842 (.ZN (CLOCK_slo__sro_n1151), .A1 (n_26), .A2 (p_0[26]));
OAI21_X2 CLOCK_slo__sro_c843 (.ZN (n_27), .A (CLOCK_slo__sro_n1152), .B1 (CLOCK_slo__sro_n1151), .B2 (CLOCK_slo__sro_n1153));
XNOR2_X2 CLOCK_slo__sro_c844 (.ZN (CLOCK_slo__sro_n1150), .A (n_26), .B (p_0[26]));
XNOR2_X1 CLOCK_slo__sro_c845 (.ZN (p_2[26]), .A (CLOCK_slo__sro_n1150), .B (p_1[26]));
INV_X1 CLOCK_slo__sro_c940 (.ZN (CLOCK_slo__sro_n1250), .A (n_15));
NAND2_X1 CLOCK_slo__sro_c941 (.ZN (CLOCK_slo__sro_n1249), .A1 (p_1[15]), .A2 (p_0[15]));
NOR2_X1 CLOCK_slo__sro_c942 (.ZN (CLOCK_slo__sro_n1248), .A1 (p_1[15]), .A2 (p_0[15]));
OAI21_X1 CLOCK_slo__sro_c943 (.ZN (CLOCK_slo__sro_n1247), .A (CLOCK_slo__sro_n1249)
    , .B1 (CLOCK_slo__sro_n1250), .B2 (CLOCK_slo__sro_n1248));
XNOR2_X1 CLOCK_slo__sro_c944 (.ZN (CLOCK_slo__sro_n1246), .A (p_1[15]), .B (p_0[15]));
XNOR2_X1 CLOCK_slo__sro_c945 (.ZN (p_2[15]), .A (CLOCK_slo__sro_n1246), .B (n_15));
OAI21_X1 CLOCK_slo__sro_c1125 (.ZN (CLOCK_slo__sro_n1442), .A (p_1[1]), .B1 (n_1), .B2 (p_0[1]));
NAND2_X1 CLOCK_slo__sro_c1126 (.ZN (n_2), .A1 (CLOCK_slo__sro_n1442), .A2 (CLOCK_slo__sro_n1443));
XNOR2_X1 CLOCK_slo__sro_c1127 (.ZN (CLOCK_slo__sro_n1441), .A (n_1), .B (p_0[1]));
XNOR2_X1 CLOCK_slo__sro_c1128 (.ZN (p_2[1]), .A (CLOCK_slo__sro_n1441), .B (p_1[1]));

endmodule //datapath__0_207

module datapath__0_206 (drc_ipoPP_0, drc_ipoPP_1, drc_ipoPP_2, Multiplier, p_0, p_1);

output [31:0] p_1;
input [31:0] Multiplier;
input [31:0] p_0;
input drc_ipoPP_0;
input drc_ipoPP_1;
input drc_ipoPP_2;
wire slo__n937;
wire n_1;
wire n_2;
wire n_3;
wire n_4;
wire n_5;
wire n_6;
wire n_7;
wire n_8;
wire n_9;
wire n_10;
wire n_11;
wire n_12;
wire n_14;
wire n_16;
wire CLOCK_slo__mro_n1915;
wire n_19;
wire n_22;
wire n_23;
wire n_24;
wire n_25;
wire n_26;
wire n_27;
wire n_29;
wire n_30;
wire n_32;
wire n_0;
wire n_34;
wire n_33;
wire slo__sro_n59;
wire slo__sro_n60;
wire slo__sro_n61;
wire slo__sro_n62;
wire slo__sro_n63;
wire slo__sro_n76;
wire slo__sro_n77;
wire slo__sro_n78;
wire slo__sro_n79;
wire slo__sro_n89;
wire slo__sro_n90;
wire slo__sro_n91;
wire slo__sro_n92;
wire slo__sro_n115;
wire slo__sro_n116;
wire slo__sro_n117;
wire slo__sro_n142;
wire slo__sro_n143;
wire slo__sro_n144;
wire slo__sro_n145;
wire slo__sro_n689;
wire slo__sro_n688;
wire slo__sro_n156;
wire slo__sro_n157;
wire slo__sro_n158;
wire slo__sro_n159;
wire slo__sro_n174;
wire slo__sro_n175;
wire slo__sro_n176;
wire slo__sro_n194;
wire slo__sro_n195;
wire slo__sro_n196;
wire slo__sro_n197;
wire slo__sro_n210;
wire slo__sro_n211;
wire slo__sro_n212;
wire slo__sro_n224;
wire CLOCK_slo__xsl_n1514;
wire slo__sro_n226;
wire slo__sro_n227;
wire slo__sro_n243;
wire slo__sro_n244;
wire slo__sro_n245;
wire slo__sro_n246;
wire slo__sro_n247;
wire slo__sro_n262;
wire slo__sro_n263;
wire slo__sro_n264;
wire slo__sro_n265;
wire slo__sro_n279;
wire slo__sro_n280;
wire slo__sro_n281;
wire slo__sro_n282;
wire slo__sro_n357;
wire slo__sro_n452;
wire slo__sro_n453;
wire slo__sro_n454;
wire slo__sro_n455;
wire slo__mro_n679;
wire slo__sro_n466;
wire slo__sro_n467;
wire slo__sro_n468;
wire slo__sro_n478;
wire slo__sro_n479;
wire slo__sro_n480;
wire slo__sro_n481;
wire slo__sro_n524;
wire slo__sro_n525;
wire slo__sro_n526;
wire slo__sro_n527;
wire slo__sro_n545;
wire slo__sro_n546;
wire slo__sro_n547;
wire slo__sro_n548;
wire slo__sro_n549;
wire slo__mro_n584;
wire slo__sro_n690;
wire slo__sro_n691;
wire slo__sro_n692;
wire slo__sro_n723;
wire slo__sro_n724;
wire slo__sro_n725;
wire slo__sro_n726;
wire slo__sro_n800;
wire slo__sro_n801;
wire slo__sro_n802;
wire slo__sro_n803;
wire slo__sro_n804;
wire slo__sro_n819;
wire slo__sro_n820;
wire slo__sro_n821;
wire slo__sro_n822;
wire slo__n940;
wire slo__sro_n943;
wire CLOCK_slo__sro_n1258;
wire CLOCK_slo__sro_n1259;
wire CLOCK_slo__sro_n1260;
wire CLOCK_slo__sro_n1261;
wire CLOCK_slo__sro_n1277;
wire CLOCK_slo__sro_n1278;
wire CLOCK_slo__sro_n1279;
wire CLOCK_slo__mro_n1326;
wire CLOCK_slo__sro_n1419;
wire CLOCK_slo__xsl_n1515;


INV_X1 i_36 (.ZN (n_34), .A (Multiplier[30]));
INV_X1 i_35 (.ZN (n_33), .A (p_0[30]));
INV_X2 i_34 (.ZN (n_32), .A (n_30));
NAND2_X1 slo__sro_c575 (.ZN (slo__sro_n726), .A1 (p_0[25]), .A2 (Multiplier[25]));
XOR2_X1 i_32 (.Z (p_1[31]), .A (slo__sro_n688), .B (Multiplier[31]));
XNOR2_X1 i_0 (.ZN (p_1[30]), .A (n_32), .B (n_0));
FA_X1 i_30 (.CO (n_30), .S (p_1[29]), .A (Multiplier[29]), .B (p_0[29]), .CI (n_29));
FA_X1 i_29 (.CO (n_29), .S (p_1[28]), .A (Multiplier[28]), .B (p_0[28]), .CI (slo__sro_n801));
INV_X1 slo__sro_c658 (.ZN (slo__sro_n822), .A (n_3));
NAND2_X1 slo__sro_c363 (.ZN (slo__sro_n481), .A1 (slo__n937), .A2 (Multiplier[17]));
INV_X1 slo__sro_c642 (.ZN (slo__sro_n804), .A (n_27));
INV_X1 slo__sro_c162 (.ZN (slo__sro_n227), .A (n_22));
INV_X1 slo__sro_c215 (.ZN (slo__sro_n282), .A (p_0[21]));
INV_X1 slo__sro_c183 (.ZN (slo__sro_n247), .A (n_19));
XNOR2_X2 slo__mro_c457 (.ZN (slo__mro_n584), .A (n_24), .B (Multiplier[24]));
INV_X1 slo__sro_c17 (.ZN (slo__sro_n79), .A (n_11));
INV_X2 slo__sro_c199 (.ZN (slo__sro_n265), .A (p_0[23]));
FA_X1 i_19 (.CO (n_19), .S (p_1[18]), .A (Multiplier[18]), .B (p_0[18]), .CI (slo__sro_n479));
INV_X1 slo__sro_c407 (.ZN (slo__sro_n527), .A (slo__sro_n546));
INV_X1 slo__sro_c132 (.ZN (slo__sro_n197), .A (n_10));
INV_X1 slo__sro_c427 (.ZN (slo__sro_n549), .A (n_14));
XNOR2_X2 slo__mro_c458 (.ZN (p_1[24]), .A (slo__mro_n584), .B (p_0[24]));
XNOR2_X2 CLOCK_slo__mro_c1697 (.ZN (CLOCK_slo__mro_n1915), .A (p_0[4]), .B (Multiplier[4]));
INV_X1 slo__sro_c113 (.ZN (slo__sro_n176), .A (n_16));
INV_X1 slo__sro_c31 (.ZN (slo__sro_n92), .A (n_6));
INV_X1 slo__sro_c146 (.ZN (slo__sro_n212), .A (n_24));
FA_X1 i_10 (.CO (n_10), .S (p_1[9]), .A (Multiplier[9]), .B (p_0[9]), .CI (n_9));
INV_X1 slo__sro_c99 (.ZN (slo__sro_n159), .A (p_0[12]));
FA_X1 i_8 (.CO (n_8), .S (p_1[7]), .A (Multiplier[7]), .B (p_0[7]), .CI (n_7));
INV_X1 slo__sro_c58 (.ZN (slo__sro_n117), .A (n_4));
XNOR2_X2 CLOCK_slo__mro_c1066 (.ZN (CLOCK_slo__mro_n1326), .A (n_26), .B (Multiplier[26]));
INV_X1 slo__sro_c85 (.ZN (slo__sro_n145), .A (n_8));
OAI21_X1 slo__c731 (.ZN (slo__n937), .A (slo__sro_n175), .B1 (slo__sro_n174), .B2 (slo__sro_n176));
FA_X1 i_3 (.CO (n_3), .S (p_1[2]), .A (Multiplier[2]), .B (p_0[2]), .CI (n_2));
INV_X1 slo__sro_c349 (.ZN (slo__sro_n468), .A (n_26));
HA_X1 i_1 (.CO (n_1), .S (p_1[0]), .A (Multiplier[0]), .B (p_0[0]));
INV_X1 slo__sro_c3 (.ZN (slo__sro_n63), .A (slo__sro_n244));
NAND2_X1 slo__sro_c4 (.ZN (slo__sro_n62), .A1 (p_0[20]), .A2 (Multiplier[20]));
NOR2_X2 slo__sro_c5 (.ZN (slo__sro_n61), .A1 (p_0[20]), .A2 (Multiplier[20]));
OAI21_X1 slo__sro_c6 (.ZN (slo__sro_n60), .A (slo__sro_n62), .B1 (slo__sro_n63), .B2 (slo__sro_n61));
XNOR2_X2 slo__sro_c7 (.ZN (slo__sro_n59), .A (p_0[20]), .B (Multiplier[20]));
XNOR2_X1 slo__sro_c8 (.ZN (p_1[20]), .A (slo__sro_n59), .B (slo__sro_n244));
NAND2_X1 slo__sro_c18 (.ZN (slo__sro_n78), .A1 (p_0[11]), .A2 (Multiplier[11]));
NOR2_X1 slo__sro_c19 (.ZN (slo__sro_n77), .A1 (p_0[11]), .A2 (Multiplier[11]));
OAI21_X2 slo__sro_c20 (.ZN (n_12), .A (slo__sro_n78), .B1 (slo__sro_n79), .B2 (slo__sro_n77));
XNOR2_X2 slo__sro_c21 (.ZN (slo__sro_n76), .A (p_0[11]), .B (Multiplier[11]));
XNOR2_X2 slo__sro_c22 (.ZN (p_1[11]), .A (slo__sro_n76), .B (n_11));
NAND2_X1 slo__sro_c32 (.ZN (slo__sro_n91), .A1 (p_0[6]), .A2 (drc_ipoPP_0));
NOR2_X1 slo__sro_c33 (.ZN (slo__sro_n90), .A1 (p_0[6]), .A2 (drc_ipoPP_0));
OAI21_X1 slo__sro_c34 (.ZN (n_7), .A (slo__sro_n91), .B1 (slo__sro_n90), .B2 (slo__sro_n92));
XNOR2_X1 slo__sro_c35 (.ZN (slo__sro_n89), .A (p_0[6]), .B (Multiplier[6]));
XNOR2_X1 slo__sro_c36 (.ZN (p_1[6]), .A (slo__sro_n89), .B (n_6));
NAND2_X1 slo__sro_c59 (.ZN (slo__sro_n116), .A1 (p_0[4]), .A2 (Multiplier[4]));
NOR2_X1 slo__sro_c60 (.ZN (slo__sro_n115), .A1 (p_0[4]), .A2 (Multiplier[4]));
OAI21_X2 slo__sro_c61 (.ZN (n_5), .A (slo__sro_n116), .B1 (slo__sro_n115), .B2 (slo__sro_n117));
OAI21_X2 CLOCK_slo__sro_c1740 (.ZN (slo__sro_n480), .A (p_0[17]), .B1 (slo__sro_n357), .B2 (Multiplier[17]));
NAND2_X1 slo__sro_c86 (.ZN (slo__sro_n144), .A1 (p_0[8]), .A2 (Multiplier[8]));
NOR2_X2 slo__sro_c87 (.ZN (slo__sro_n143), .A1 (p_0[8]), .A2 (drc_ipoPP_1));
OAI21_X2 slo__sro_c88 (.ZN (n_9), .A (slo__sro_n144), .B1 (slo__sro_n143), .B2 (slo__sro_n145));
XNOR2_X1 slo__sro_c89 (.ZN (slo__sro_n142), .A (p_0[8]), .B (Multiplier[8]));
XNOR2_X1 slo__sro_c90 (.ZN (p_1[8]), .A (slo__sro_n142), .B (n_8));
NAND2_X1 slo__sro_c100 (.ZN (slo__sro_n158), .A1 (n_12), .A2 (Multiplier[12]));
NOR2_X1 slo__sro_c101 (.ZN (slo__sro_n157), .A1 (n_12), .A2 (Multiplier[12]));
OAI21_X1 slo__sro_c102 (.ZN (slo__sro_n156), .A (slo__sro_n158), .B1 (slo__sro_n159), .B2 (slo__sro_n157));
INV_X1 slo__sro_c544 (.ZN (slo__sro_n692), .A (n_30));
NOR2_X1 slo__sro_c545 (.ZN (slo__sro_n691), .A1 (n_33), .A2 (Multiplier[30]));
NAND2_X1 slo__sro_c114 (.ZN (slo__sro_n175), .A1 (p_0[16]), .A2 (Multiplier[16]));
NOR2_X2 slo__sro_c115 (.ZN (slo__sro_n174), .A1 (p_0[16]), .A2 (Multiplier[16]));
INV_X1 slo__sro_c335 (.ZN (slo__sro_n455), .A (p_0[1]));
INV_X1 CLOCK_slo__sro_c999 (.ZN (CLOCK_slo__sro_n1261), .A (slo__sro_n156));
XNOR2_X1 slo__sro_c118 (.ZN (p_1[16]), .A (slo__sro_n943), .B (n_16));
NAND2_X1 slo__sro_c133 (.ZN (slo__sro_n196), .A1 (p_0[10]), .A2 (Multiplier[10]));
NOR2_X1 slo__sro_c134 (.ZN (slo__sro_n195), .A1 (p_0[10]), .A2 (Multiplier[10]));
OAI21_X2 slo__sro_c135 (.ZN (n_11), .A (slo__sro_n196), .B1 (slo__sro_n197), .B2 (slo__sro_n195));
XNOR2_X1 slo__sro_c136 (.ZN (slo__sro_n194), .A (p_0[10]), .B (Multiplier[10]));
NAND2_X1 slo__sro_c147 (.ZN (slo__sro_n211), .A1 (p_0[24]), .A2 (Multiplier[24]));
NOR2_X1 CLOCK_slo__sro_c1001 (.ZN (CLOCK_slo__sro_n1259), .A1 (p_0[13]), .A2 (Multiplier[13]));
OAI21_X2 slo__sro_c149 (.ZN (n_25), .A (slo__sro_n211), .B1 (slo__sro_n210), .B2 (slo__sro_n212));
XNOR2_X1 slo__mro_c513 (.ZN (p_1[10]), .A (n_10), .B (slo__sro_n194));
OAI22_X1 CLOCK_slo__sro_c1235 (.ZN (n_0), .A1 (n_33), .A2 (Multiplier[30]), .B1 (p_0[30]), .B2 (n_34));
NAND2_X2 slo__sro_c163 (.ZN (slo__sro_n226), .A1 (p_0[22]), .A2 (Multiplier[22]));
INV_X1 CLOCK_slo__xsl_c1260 (.ZN (CLOCK_slo__xsl_n1514), .A (CLOCK_slo__xsl_n1515));
OAI21_X2 slo__sro_c165 (.ZN (n_23), .A (slo__sro_n226), .B1 (CLOCK_slo__sro_n1419), .B2 (slo__sro_n227));
XNOR2_X1 slo__sro_c166 (.ZN (slo__sro_n224), .A (p_0[22]), .B (Multiplier[22]));
XNOR2_X2 slo__sro_c167 (.ZN (p_1[22]), .A (slo__sro_n224), .B (n_22));
NAND2_X1 slo__sro_c184 (.ZN (slo__sro_n246), .A1 (p_0[19]), .A2 (Multiplier[19]));
NOR2_X1 slo__sro_c185 (.ZN (slo__sro_n245), .A1 (p_0[19]), .A2 (Multiplier[19]));
OAI21_X2 slo__sro_c186 (.ZN (slo__sro_n244), .A (slo__sro_n246), .B1 (slo__sro_n247), .B2 (slo__sro_n245));
XNOR2_X2 slo__sro_c187 (.ZN (slo__sro_n243), .A (p_0[19]), .B (Multiplier[19]));
XNOR2_X2 slo__sro_c188 (.ZN (p_1[19]), .A (n_19), .B (slo__sro_n243));
NAND2_X1 slo__sro_c200 (.ZN (slo__sro_n264), .A1 (n_23), .A2 (Multiplier[23]));
NOR2_X1 slo__sro_c201 (.ZN (slo__sro_n263), .A1 (n_23), .A2 (Multiplier[23]));
OAI21_X2 slo__sro_c202 (.ZN (n_24), .A (slo__sro_n264), .B1 (slo__sro_n265), .B2 (slo__sro_n263));
XNOR2_X2 slo__sro_c203 (.ZN (slo__sro_n262), .A (n_23), .B (Multiplier[23]));
XNOR2_X1 slo__sro_c204 (.ZN (p_1[23]), .A (slo__sro_n262), .B (p_0[23]));
NAND2_X1 slo__sro_c216 (.ZN (slo__sro_n281), .A1 (slo__sro_n60), .A2 (Multiplier[21]));
NOR2_X1 slo__sro_c217 (.ZN (slo__sro_n280), .A1 (slo__sro_n60), .A2 (Multiplier[21]));
OAI21_X2 slo__sro_c218 (.ZN (n_22), .A (slo__sro_n281), .B1 (slo__sro_n280), .B2 (slo__sro_n282));
XNOR2_X1 slo__sro_c219 (.ZN (slo__sro_n279), .A (slo__n940), .B (Multiplier[21]));
XNOR2_X1 slo__sro_c220 (.ZN (p_1[21]), .A (slo__sro_n279), .B (p_0[21]));
OAI21_X2 slo__sro_c275 (.ZN (slo__sro_n357), .A (slo__sro_n175), .B1 (slo__sro_n174), .B2 (slo__sro_n176));
NAND2_X1 slo__sro_c336 (.ZN (slo__sro_n454), .A1 (n_1), .A2 (Multiplier[1]));
NOR2_X1 slo__sro_c337 (.ZN (slo__sro_n453), .A1 (n_1), .A2 (Multiplier[1]));
OAI21_X1 slo__sro_c338 (.ZN (n_2), .A (slo__sro_n454), .B1 (slo__sro_n455), .B2 (slo__sro_n453));
XNOR2_X1 slo__sro_c339 (.ZN (slo__sro_n452), .A (n_1), .B (Multiplier[1]));
XNOR2_X1 slo__sro_c340 (.ZN (p_1[1]), .A (slo__sro_n452), .B (p_0[1]));
NAND2_X1 slo__sro_c350 (.ZN (slo__sro_n467), .A1 (p_0[26]), .A2 (Multiplier[26]));
NOR2_X1 slo__sro_c351 (.ZN (slo__sro_n466), .A1 (p_0[26]), .A2 (Multiplier[26]));
OAI21_X2 slo__sro_c352 (.ZN (n_27), .A (slo__sro_n467), .B1 (slo__sro_n466), .B2 (slo__sro_n468));
XNOR2_X1 slo__mro_c536 (.ZN (slo__mro_n679), .A (p_0[12]), .B (Multiplier[12]));
XNOR2_X1 slo__mro_c537 (.ZN (p_1[12]), .A (slo__mro_n679), .B (n_12));
NAND2_X2 slo__sro_c365 (.ZN (slo__sro_n479), .A1 (slo__sro_n480), .A2 (slo__sro_n481));
XNOR2_X1 slo__sro_c366 (.ZN (slo__sro_n478), .A (p_0[17]), .B (Multiplier[17]));
XNOR2_X1 slo__sro_c367 (.ZN (p_1[17]), .A (slo__sro_n478), .B (slo__sro_n357));
NAND2_X1 slo__sro_c408 (.ZN (slo__sro_n526), .A1 (p_0[15]), .A2 (Multiplier[15]));
NOR2_X1 slo__sro_c409 (.ZN (slo__sro_n525), .A1 (p_0[15]), .A2 (Multiplier[15]));
OAI21_X2 slo__sro_c410 (.ZN (n_16), .A (slo__sro_n526), .B1 (slo__sro_n527), .B2 (slo__sro_n525));
XNOR2_X2 slo__sro_c411 (.ZN (slo__sro_n524), .A (p_0[15]), .B (Multiplier[15]));
XNOR2_X2 slo__sro_c412 (.ZN (p_1[15]), .A (slo__sro_n524), .B (slo__sro_n546));
NAND2_X1 slo__sro_c428 (.ZN (slo__sro_n548), .A1 (p_0[14]), .A2 (Multiplier[14]));
NOR2_X1 slo__sro_c429 (.ZN (slo__sro_n547), .A1 (p_0[14]), .A2 (Multiplier[14]));
OAI21_X2 slo__sro_c430 (.ZN (slo__sro_n546), .A (slo__sro_n548), .B1 (slo__sro_n547), .B2 (slo__sro_n549));
XNOR2_X1 slo__sro_c431 (.ZN (slo__sro_n545), .A (p_0[14]), .B (Multiplier[14]));
XNOR2_X1 slo__sro_c432 (.ZN (p_1[14]), .A (slo__sro_n545), .B (n_14));
NAND2_X1 slo__sro_c546 (.ZN (slo__sro_n690), .A1 (slo__sro_n692), .A2 (slo__sro_n691));
OR2_X1 slo__sro_c547 (.ZN (slo__sro_n689), .A1 (p_0[30]), .A2 (n_34));
OAI21_X1 slo__sro_c548 (.ZN (slo__sro_n688), .A (slo__sro_n690), .B1 (n_32), .B2 (slo__sro_n689));
NAND2_X2 slo__sro_c576 (.ZN (slo__sro_n725), .A1 (n_25), .A2 (Multiplier[25]));
NAND2_X2 slo__sro_c577 (.ZN (slo__sro_n724), .A1 (n_25), .A2 (p_0[25]));
NAND3_X2 slo__sro_c578 (.ZN (n_26), .A1 (slo__sro_n725), .A2 (slo__sro_n724), .A3 (slo__sro_n726));
XNOR2_X1 slo__sro_c579 (.ZN (slo__sro_n723), .A (p_0[25]), .B (Multiplier[25]));
XNOR2_X1 slo__sro_c580 (.ZN (p_1[25]), .A (slo__sro_n723), .B (n_25));
NAND2_X1 slo__sro_c643 (.ZN (slo__sro_n803), .A1 (p_0[27]), .A2 (Multiplier[27]));
NOR2_X2 slo__sro_c644 (.ZN (slo__sro_n802), .A1 (p_0[27]), .A2 (Multiplier[27]));
OAI21_X1 slo__sro_c645 (.ZN (slo__sro_n801), .A (slo__sro_n803), .B1 (slo__sro_n804), .B2 (slo__sro_n802));
XNOR2_X2 slo__sro_c646 (.ZN (slo__sro_n800), .A (p_0[27]), .B (Multiplier[27]));
XNOR2_X1 slo__sro_c647 (.ZN (p_1[27]), .A (slo__sro_n800), .B (n_27));
NAND2_X1 slo__sro_c659 (.ZN (slo__sro_n821), .A1 (p_0[3]), .A2 (Multiplier[3]));
NOR2_X1 slo__sro_c660 (.ZN (slo__sro_n820), .A1 (p_0[3]), .A2 (Multiplier[3]));
OAI21_X2 slo__sro_c661 (.ZN (n_4), .A (slo__sro_n821), .B1 (slo__sro_n822), .B2 (slo__sro_n820));
XNOR2_X2 slo__sro_c662 (.ZN (slo__sro_n819), .A (p_0[3]), .B (Multiplier[3]));
XNOR2_X1 slo__sro_c663 (.ZN (p_1[3]), .A (slo__sro_n819), .B (n_3));
OAI21_X1 slo__c734 (.ZN (slo__n940), .A (slo__sro_n62), .B1 (slo__sro_n63), .B2 (slo__sro_n61));
XNOR2_X1 slo__sro_c737 (.ZN (slo__sro_n943), .A (p_0[16]), .B (drc_ipoPP_2));
NAND2_X1 CLOCK_slo__sro_c1000 (.ZN (CLOCK_slo__sro_n1260), .A1 (p_0[13]), .A2 (Multiplier[13]));
NOR2_X2 CLOCK_slo__mro_c986 (.ZN (slo__sro_n210), .A1 (p_0[24]), .A2 (Multiplier[24]));
OAI21_X1 CLOCK_slo__sro_c1002 (.ZN (n_14), .A (CLOCK_slo__sro_n1260), .B1 (CLOCK_slo__sro_n1259), .B2 (CLOCK_slo__sro_n1261));
XNOR2_X2 CLOCK_slo__sro_c1003 (.ZN (CLOCK_slo__sro_n1258), .A (p_0[13]), .B (Multiplier[13]));
XNOR2_X2 CLOCK_slo__sro_c1004 (.ZN (p_1[13]), .A (CLOCK_slo__sro_n1258), .B (CLOCK_slo__xsl_n1514));
NAND2_X1 CLOCK_slo__sro_c1021 (.ZN (CLOCK_slo__sro_n1279), .A1 (p_0[5]), .A2 (Multiplier[5]));
AOI22_X1 CLOCK_slo__sro_c1022 (.ZN (CLOCK_slo__sro_n1278), .A1 (p_0[5]), .A2 (n_5)
    , .B1 (n_5), .B2 (Multiplier[5]));
NAND2_X1 CLOCK_slo__sro_c1023 (.ZN (n_6), .A1 (CLOCK_slo__sro_n1278), .A2 (CLOCK_slo__sro_n1279));
XNOR2_X1 CLOCK_slo__sro_c1024 (.ZN (CLOCK_slo__sro_n1277), .A (n_5), .B (Multiplier[5]));
XNOR2_X1 CLOCK_slo__sro_c1025 (.ZN (p_1[5]), .A (CLOCK_slo__sro_n1277), .B (p_0[5]));
XNOR2_X2 CLOCK_slo__mro_c1067 (.ZN (p_1[26]), .A (CLOCK_slo__mro_n1326), .B (p_0[26]));
INV_X1 CLOCK_slo__xsl_c1259 (.ZN (CLOCK_slo__xsl_n1515), .A (slo__sro_n156));
NOR2_X2 CLOCK_slo__sro_c1175 (.ZN (CLOCK_slo__sro_n1419), .A1 (p_0[22]), .A2 (Multiplier[22]));
XNOR2_X2 CLOCK_slo__mro_c1698 (.ZN (p_1[4]), .A (CLOCK_slo__mro_n1915), .B (n_4));

endmodule //datapath__0_206

module datapath__0_202 (p_0, p_1, p_2);

output [31:0] p_2;
input [31:0] p_0;
input [31:0] p_1;
wire CLOCK_slo__mro_n1501;
wire slo__sro_n601;
wire n_1;
wire n_2;
wire n_3;
wire n_4;
wire n_5;
wire n_6;
wire n_7;
wire n_8;
wire n_9;
wire n_10;
wire n_11;
wire n_12;
wire n_13;
wire n_14;
wire n_16;
wire n_17;
wire n_18;
wire n_19;
wire n_20;
wire n_22;
wire n_25;
wire n_26;
wire n_27;
wire n_28;
wire n_29;
wire n_30;
wire n_32;
wire n_0;
wire n_34;
wire n_33;
wire n_31;
wire slo__sro_n63;
wire slo__sro_n64;
wire slo__sro_n65;
wire slo__sro_n66;
wire slo__sro_n78;
wire slo__sro_n79;
wire slo__sro_n80;
wire slo__sro_n81;
wire slo__sro_n93;
wire slo__sro_n94;
wire slo__sro_n95;
wire slo__sro_n96;
wire slo__sro_n121;
wire slo__sro_n122;
wire slo__sro_n123;
wire slo__sro_n124;
wire slo__sro_n125;
wire slo__sro_n138;
wire slo__sro_n139;
wire slo__sro_n141;
wire slo__sro_n167;
wire slo__sro_n168;
wire slo__sro_n169;
wire slo__sro_n170;
wire slo__sro_n171;
wire slo__sro_n172;
wire slo__sro_n184;
wire slo__sro_n185;
wire slo__sro_n186;
wire slo__sro_n187;
wire slo__sro_n286;
wire slo__sro_n287;
wire slo__sro_n288;
wire slo__sro_n289;
wire slo__sro_n452;
wire slo__sro_n453;
wire slo__sro_n454;
wire slo__sro_n544;
wire slo__sro_n545;
wire slo__n820;
wire slo__sro_n547;
wire slo__sro_n602;
wire slo__sro_n603;
wire CLOCK_sgo__sro_n958;
wire CLOCK_sgo__sro_n959;
wire CLOCK_sgo__sro_n960;
wire CLOCK_sgo__sro_n961;
wire CLOCK_slo__sro_n1015;
wire CLOCK_slo__sro_n1016;
wire CLOCK_slo__sro_n1017;
wire CLOCK_slo__sro_n1018;
wire CLOCK_slo__sro_n1074;
wire CLOCK_slo__sro_n1075;
wire CLOCK_slo__sro_n1076;
wire CLOCK_slo__sro_n1077;
wire CLOCK_slo__sro_n1078;
wire CLOCK_slo__sro_n1150;
wire CLOCK_slo__sro_n1151;
wire CLOCK_slo__sro_n1152;
wire CLOCK_slo__sro_n1414;
wire CLOCK_slo__sro_n1415;
wire CLOCK_slo__sro_n1416;
wire CLOCK_slo__sro_n1118;
wire CLOCK_slo__sro_n1119;
wire CLOCK_slo__sro_n1120;
wire CLOCK_slo__sro_n1121;


INV_X1 i_36 (.ZN (n_34), .A (p_0[30]));
INV_X1 i_35 (.ZN (n_33), .A (p_1[30]));
INV_X1 i_34 (.ZN (n_32), .A (n_30));
XNOR2_X2 CLOCK_slo__mro_c1075 (.ZN (CLOCK_slo__mro_n1501), .A (p_1[25]), .B (p_0[25]));
XOR2_X1 i_32 (.Z (p_2[31]), .A (p_0[31]), .B (n_31));
OAI22_X1 i_31 (.ZN (n_0), .A1 (n_34), .A2 (p_1[30]), .B1 (p_0[30]), .B2 (n_33));
XNOR2_X1 i_0 (.ZN (p_2[30]), .A (n_32), .B (n_0));
FA_X1 i_30 (.CO (n_30), .S (p_2[29]), .A (p_0[29]), .B (p_1[29]), .CI (n_29));
FA_X1 i_28 (.CO (n_28), .S (p_2[27]), .A (p_0[27]), .B (p_1[27]), .CI (n_27));
NAND2_X1 slo__sro_c324 (.ZN (slo__sro_n547), .A1 (p_0[23]), .A2 (p_1[23]));
FA_X1 i_25 (.CO (n_25), .S (p_2[24]), .A (p_0[24]), .B (p_1[24]), .CI (slo__sro_n545));
NOR2_X1 slo__sro_c357 (.ZN (slo__sro_n603), .A1 (p_1[23]), .A2 (p_0[23]));
INV_X1 slo__sro_c99 (.ZN (slo__sro_n172), .A (p_0[1]));
FA_X1 i_22 (.CO (n_22), .S (p_2[21]), .A (p_0[21]), .B (p_1[21]), .CI (slo__sro_n122));
NAND2_X1 slo__sro_c72 (.ZN (slo__sro_n141), .A1 (p_1[22]), .A2 (p_0[22]));
INV_X2 slo__sro_c17 (.ZN (slo__sro_n81), .A (n_18));
INV_X2 slo__sro_c31 (.ZN (slo__sro_n96), .A (n_11));
FA_X1 i_18 (.CO (n_18), .S (p_2[17]), .A (p_0[17]), .B (p_1[17]), .CI (n_17));
FA_X1 i_17 (.CO (n_17), .S (p_2[16]), .A (p_0[16]), .B (p_1[16]), .CI (n_16));
FA_X1 i_16 (.CO (n_16), .S (p_2[15]), .A (p_0[15]), .B (p_1[15]), .CI (CLOCK_slo__sro_n1075));
NAND2_X1 CLOCK_slo__sro_c795 (.ZN (CLOCK_slo__sro_n1152), .A1 (p_1[28]), .A2 (p_0[28]));
FA_X1 i_14 (.CO (n_14), .S (p_2[13]), .A (p_0[13]), .B (p_1[13]), .CI (n_13));
INV_X1 slo__sro_c169 (.ZN (slo__sro_n289), .A (n_30));
INV_X1 slo__sro_c58 (.ZN (slo__sro_n125), .A (n_20));
INV_X1 CLOCK_slo__sro_c720 (.ZN (CLOCK_slo__sro_n1078), .A (n_14));
FA_X1 i_10 (.CO (n_10), .S (p_2[9]), .A (p_0[9]), .B (p_1[9]), .CI (n_9));
FA_X1 i_9 (.CO (n_9), .S (p_2[8]), .A (p_0[8]), .B (p_1[8]), .CI (n_8));
FA_X1 i_8 (.CO (n_8), .S (p_2[7]), .A (p_0[7]), .B (p_1[7]), .CI (n_7));
FA_X1 i_7 (.CO (n_7), .S (p_2[6]), .A (p_0[6]), .B (p_1[6]), .CI (n_6));
FA_X1 i_5 (.CO (n_5), .S (p_2[4]), .A (p_0[4]), .B (p_1[4]), .CI (n_4));
FA_X1 i_4 (.CO (n_4), .S (p_2[3]), .A (p_0[3]), .B (p_1[3]), .CI (n_3));
FA_X1 i_3 (.CO (n_3), .S (p_2[2]), .A (p_0[2]), .B (p_1[2]), .CI (n_2));
INV_X1 slo__sro_c117 (.ZN (slo__sro_n187), .A (n_12));
HA_X1 i_1 (.CO (n_1), .S (p_2[0]), .A (p_0[0]), .B (p_1[0]));
INV_X2 slo__sro_c1 (.ZN (slo__sro_n66), .A (slo__n820));
NAND2_X1 slo__sro_c2 (.ZN (slo__sro_n65), .A1 (p_1[19]), .A2 (p_0[19]));
NOR2_X1 slo__sro_c3 (.ZN (slo__sro_n64), .A1 (p_1[19]), .A2 (p_0[19]));
OAI21_X2 slo__sro_c4 (.ZN (n_20), .A (slo__sro_n65), .B1 (slo__sro_n64), .B2 (slo__sro_n66));
XNOR2_X1 slo__sro_c5 (.ZN (slo__sro_n63), .A (p_1[19]), .B (p_0[19]));
XNOR2_X2 slo__sro_c6 (.ZN (p_2[19]), .A (n_19), .B (slo__sro_n63));
NAND2_X1 slo__sro_c18 (.ZN (slo__sro_n80), .A1 (p_1[18]), .A2 (p_0[18]));
NOR2_X1 slo__sro_c19 (.ZN (slo__sro_n79), .A1 (p_1[18]), .A2 (p_0[18]));
OAI21_X2 slo__sro_c20 (.ZN (n_19), .A (slo__sro_n80), .B1 (slo__sro_n81), .B2 (slo__sro_n79));
XNOR2_X1 slo__sro_c21 (.ZN (slo__sro_n78), .A (p_1[18]), .B (p_0[18]));
XNOR2_X1 slo__sro_c22 (.ZN (p_2[18]), .A (n_18), .B (slo__sro_n78));
NAND2_X1 slo__sro_c32 (.ZN (slo__sro_n95), .A1 (p_1[11]), .A2 (p_0[11]));
NOR2_X1 slo__sro_c33 (.ZN (slo__sro_n94), .A1 (p_1[11]), .A2 (p_0[11]));
OAI21_X2 slo__sro_c34 (.ZN (n_12), .A (slo__sro_n95), .B1 (slo__sro_n96), .B2 (slo__sro_n94));
XNOR2_X1 slo__sro_c35 (.ZN (slo__sro_n93), .A (p_1[11]), .B (p_0[11]));
XNOR2_X1 slo__sro_c36 (.ZN (p_2[11]), .A (slo__sro_n93), .B (n_11));
NAND2_X1 slo__sro_c59 (.ZN (slo__sro_n124), .A1 (p_1[20]), .A2 (p_0[20]));
NOR2_X1 slo__sro_c60 (.ZN (slo__sro_n123), .A1 (p_1[20]), .A2 (p_0[20]));
OAI21_X1 slo__sro_c61 (.ZN (slo__sro_n122), .A (slo__sro_n124), .B1 (slo__sro_n125), .B2 (slo__sro_n123));
XNOR2_X1 slo__sro_c62 (.ZN (slo__sro_n121), .A (p_1[20]), .B (p_0[20]));
XNOR2_X1 slo__sro_c63 (.ZN (p_2[20]), .A (slo__sro_n121), .B (n_20));
INV_X2 CLOCK_slo__sro_c658 (.ZN (CLOCK_slo__sro_n1018), .A (n_10));
NAND2_X1 slo__sro_c74 (.ZN (slo__sro_n139), .A1 (CLOCK_sgo__sro_n958), .A2 (slo__sro_n141));
XNOR2_X1 slo__sro_c75 (.ZN (slo__sro_n138), .A (n_22), .B (p_0[22]));
XNOR2_X1 slo__sro_c76 (.ZN (p_2[22]), .A (slo__sro_n138), .B (p_1[22]));
INV_X1 slo__sro_c100 (.ZN (slo__sro_n171), .A (n_1));
NAND2_X1 slo__sro_c101 (.ZN (slo__sro_n170), .A1 (n_1), .A2 (p_0[1]));
NAND2_X1 slo__sro_c102 (.ZN (slo__sro_n169), .A1 (slo__sro_n171), .A2 (slo__sro_n172));
NAND2_X1 slo__sro_c103 (.ZN (slo__sro_n168), .A1 (p_1[1]), .A2 (slo__sro_n169));
NAND2_X1 slo__sro_c104 (.ZN (n_2), .A1 (slo__sro_n168), .A2 (slo__sro_n170));
XNOR2_X1 slo__sro_c105 (.ZN (slo__sro_n167), .A (n_1), .B (p_0[1]));
XNOR2_X1 slo__sro_c106 (.ZN (p_2[1]), .A (p_1[1]), .B (slo__sro_n167));
NAND2_X1 slo__sro_c118 (.ZN (slo__sro_n186), .A1 (p_1[12]), .A2 (p_0[12]));
NOR2_X1 slo__sro_c119 (.ZN (slo__sro_n185), .A1 (p_1[12]), .A2 (p_0[12]));
OAI21_X1 slo__sro_c120 (.ZN (n_13), .A (slo__sro_n186), .B1 (slo__sro_n187), .B2 (slo__sro_n185));
XNOR2_X1 slo__sro_c121 (.ZN (slo__sro_n184), .A (p_1[12]), .B (p_0[12]));
XNOR2_X1 slo__sro_c122 (.ZN (p_2[12]), .A (slo__sro_n184), .B (n_12));
NOR2_X1 slo__sro_c170 (.ZN (slo__sro_n288), .A1 (n_33), .A2 (p_0[30]));
NAND2_X1 slo__sro_c171 (.ZN (slo__sro_n287), .A1 (slo__sro_n288), .A2 (slo__sro_n289));
OR2_X1 slo__sro_c172 (.ZN (slo__sro_n286), .A1 (p_1[30]), .A2 (n_34));
OAI21_X1 slo__sro_c173 (.ZN (n_31), .A (slo__sro_n287), .B1 (n_32), .B2 (slo__sro_n286));
XNOR2_X2 CLOCK_slo__mro_c1076 (.ZN (p_2[25]), .A (CLOCK_slo__mro_n1501), .B (n_25));
INV_X1 slo__sro_c253 (.ZN (slo__sro_n454), .A (n_25));
NAND2_X1 slo__sro_c254 (.ZN (slo__sro_n453), .A1 (p_1[25]), .A2 (p_0[25]));
NOR2_X1 slo__sro_c255 (.ZN (slo__sro_n452), .A1 (p_1[25]), .A2 (p_0[25]));
OAI21_X1 slo__sro_c256 (.ZN (n_26), .A (slo__sro_n453), .B1 (slo__sro_n454), .B2 (slo__sro_n452));
OAI21_X1 slo__c486 (.ZN (slo__n820), .A (slo__sro_n80), .B1 (slo__sro_n81), .B2 (slo__sro_n79));
NAND2_X1 slo__sro_c326 (.ZN (slo__sro_n545), .A1 (slo__sro_n547), .A2 (slo__sro_n601));
XNOR2_X1 slo__sro_c327 (.ZN (slo__sro_n544), .A (p_1[23]), .B (p_0[23]));
XNOR2_X1 slo__sro_c328 (.ZN (p_2[23]), .A (slo__sro_n544), .B (slo__sro_n139));
INV_X1 slo__sro_c358 (.ZN (slo__sro_n602), .A (slo__sro_n603));
NAND2_X1 slo__sro_c359 (.ZN (slo__sro_n601), .A1 (slo__sro_n139), .A2 (slo__sro_n602));
INV_X1 CLOCK_sgo__sro_c589 (.ZN (CLOCK_sgo__sro_n961), .A (p_1[22]));
INV_X1 CLOCK_sgo__sro_c590 (.ZN (CLOCK_sgo__sro_n960), .A (p_0[22]));
NAND2_X1 CLOCK_sgo__sro_c591 (.ZN (CLOCK_sgo__sro_n959), .A1 (CLOCK_sgo__sro_n960), .A2 (CLOCK_sgo__sro_n961));
NAND2_X1 CLOCK_sgo__sro_c592 (.ZN (CLOCK_sgo__sro_n958), .A1 (n_22), .A2 (CLOCK_sgo__sro_n959));
NAND2_X1 CLOCK_slo__sro_c659 (.ZN (CLOCK_slo__sro_n1017), .A1 (p_1[10]), .A2 (p_0[10]));
NOR2_X1 CLOCK_slo__sro_c660 (.ZN (CLOCK_slo__sro_n1016), .A1 (p_1[10]), .A2 (p_0[10]));
OAI21_X2 CLOCK_slo__sro_c661 (.ZN (n_11), .A (CLOCK_slo__sro_n1017), .B1 (CLOCK_slo__sro_n1018), .B2 (CLOCK_slo__sro_n1016));
XNOR2_X1 CLOCK_slo__sro_c662 (.ZN (CLOCK_slo__sro_n1015), .A (p_1[10]), .B (p_0[10]));
XNOR2_X1 CLOCK_slo__sro_c663 (.ZN (p_2[10]), .A (CLOCK_slo__sro_n1015), .B (n_10));
NAND2_X1 CLOCK_slo__sro_c721 (.ZN (CLOCK_slo__sro_n1077), .A1 (p_1[14]), .A2 (p_0[14]));
NOR2_X1 CLOCK_slo__sro_c722 (.ZN (CLOCK_slo__sro_n1076), .A1 (p_1[14]), .A2 (p_0[14]));
OAI21_X1 CLOCK_slo__sro_c723 (.ZN (CLOCK_slo__sro_n1075), .A (CLOCK_slo__sro_n1077)
    , .B1 (CLOCK_slo__sro_n1078), .B2 (CLOCK_slo__sro_n1076));
XNOR2_X1 CLOCK_slo__sro_c724 (.ZN (CLOCK_slo__sro_n1074), .A (p_1[14]), .B (p_0[14]));
XNOR2_X1 CLOCK_slo__sro_c725 (.ZN (p_2[14]), .A (CLOCK_slo__sro_n1074), .B (n_14));
OAI21_X1 CLOCK_slo__sro_c796 (.ZN (CLOCK_slo__sro_n1151), .A (n_28), .B1 (p_1[28]), .B2 (p_0[28]));
NAND2_X2 CLOCK_slo__sro_c797 (.ZN (n_29), .A1 (CLOCK_slo__sro_n1151), .A2 (CLOCK_slo__sro_n1152));
XNOR2_X1 CLOCK_slo__sro_c798 (.ZN (CLOCK_slo__sro_n1150), .A (p_1[28]), .B (p_0[28]));
XNOR2_X1 CLOCK_slo__sro_c799 (.ZN (p_2[28]), .A (CLOCK_slo__sro_n1150), .B (n_28));
NAND2_X1 CLOCK_slo__sro_c990 (.ZN (CLOCK_slo__sro_n1416), .A1 (p_1[26]), .A2 (p_0[26]));
OAI21_X1 CLOCK_slo__sro_c991 (.ZN (CLOCK_slo__sro_n1415), .A (n_26), .B1 (p_1[26]), .B2 (p_0[26]));
NAND2_X1 CLOCK_slo__sro_c992 (.ZN (n_27), .A1 (CLOCK_slo__sro_n1415), .A2 (CLOCK_slo__sro_n1416));
XNOR2_X1 CLOCK_slo__sro_c993 (.ZN (CLOCK_slo__sro_n1414), .A (p_1[26]), .B (p_0[26]));
XNOR2_X1 CLOCK_slo__sro_c994 (.ZN (p_2[26]), .A (CLOCK_slo__sro_n1414), .B (n_26));
INV_X2 CLOCK_slo__sro_c762 (.ZN (CLOCK_slo__sro_n1121), .A (n_5));
NAND2_X1 CLOCK_slo__sro_c763 (.ZN (CLOCK_slo__sro_n1120), .A1 (p_1[5]), .A2 (p_0[5]));
NOR2_X1 CLOCK_slo__sro_c764 (.ZN (CLOCK_slo__sro_n1119), .A1 (p_1[5]), .A2 (p_0[5]));
OAI21_X2 CLOCK_slo__sro_c765 (.ZN (n_6), .A (CLOCK_slo__sro_n1120), .B1 (CLOCK_slo__sro_n1121), .B2 (CLOCK_slo__sro_n1119));
XNOR2_X1 CLOCK_slo__sro_c766 (.ZN (CLOCK_slo__sro_n1118), .A (p_1[5]), .B (p_0[5]));
XNOR2_X1 CLOCK_slo__sro_c767 (.ZN (p_2[5]), .A (CLOCK_slo__sro_n1118), .B (n_5));

endmodule //datapath__0_202

module datapath__0_201 (p_0_17_PP_1, opt_ipoPP_0, p_0_16_PP_5, Multiplier, p_0, p_1);

output [31:0] p_1;
input [31:0] Multiplier;
input [31:0] p_0;
input p_0_17_PP_1;
input opt_ipoPP_0;
input p_0_16_PP_5;
wire slo_n951;
wire CLOCK_slo__sro_n1695;
wire CLOCK_slo__sro_n1807;
wire slo__mro_n724;
wire CLOCK_slo__sro_n1872;
wire n_1;
wire n_2;
wire n_3;
wire slo__sro_n886;
wire n_7;
wire n_8;
wire n_9;
wire n_10;
wire n_11;
wire n_14;
wire n_15;
wire n_16;
wire n_19;
wire n_20;
wire n_21;
wire n_22;
wire n_23;
wire n_24;
wire n_25;
wire n_26;
wire n_27;
wire n_28;
wire n_30;
wire n_32;
wire n_0;
wire n_34;
wire n_33;
wire n_31;
wire slo__sro_n847;
wire slo__sro_n846;
wire slo__sro_n60;
wire slo__sro_n61;
wire slo__sro_n62;
wire slo__sro_n750;
wire slo__sro_n73;
wire slo__sro_n74;
wire slo__sro_n75;
wire slo__sro_n85;
wire slo__sro_n87;
wire slo__sro_n88;
wire slo__sro_n98;
wire slo__sro_n99;
wire slo__sro_n100;
wire slo__sro_n101;
wire slo__sro_n102;
wire slo__sro_n167;
wire slo__sro_n168;
wire slo__sro_n169;
wire slo__sro_n170;
wire slo__sro_n171;
wire slo__sro_n185;
wire slo__sro_n187;
wire slo__sro_n188;
wire slo__sro_n228;
wire slo__sro_n229;
wire slo__sro_n230;
wire slo__sro_n231;
wire slo__sro_n245;
wire slo__sro_n246;
wire slo__sro_n247;
wire slo__sro_n248;
wire slo__sro_n249;
wire slo__sro_n262;
wire slo__sro_n263;
wire slo__sro_n832;
wire slo__sro_n265;
wire slo__sro_n280;
wire slo__sro_n281;
wire slo__sro_n282;
wire slo__sro_n283;
wire CLOCK_slo__sro_n1464;
wire slo__sro_n299;
wire slo__sro_n751;
wire slo__sro_n752;
wire slo__sro_n753;
wire slo__mro_n826;
wire slo__sro_n833;
wire slo__sro_n834;
wire slo__sro_n845;
wire slo__mro_n796;
wire slo__sro_n848;
wire slo__mro_n875;
wire slo__sro_n887;
wire slo__sro_n888;
wire slo__sro_n990;
wire slo__sro_n991;
wire slo__sro_n992;
wire slo__sro_n993;
wire slo__sro_n1234;
wire CLOCK_slo__sro_n1419;
wire CLOCK_slo__sro_n1420;
wire CLOCK_slo__sro_n1421;
wire CLOCK_slo__sro_n1422;
wire CLOCK_slo__mro_n1455;
wire CLOCK_slo__sro_n1694;
wire CLOCK_slo__sro_n1486;
wire CLOCK_slo__sro_n1487;
wire CLOCK_slo__sro_n1488;
wire CLOCK_slo__sro_n1489;
wire CLOCK_slo__sro_n1696;
wire CLOCK_slo__sro_n1808;
wire CLOCK_slo__sro_n1809;
wire CLOCK_slo__sro_n1810;
wire CLOCK_slo__sro_n1873;
wire CLOCK_slo__sro_n1874;
wire CLOCK_slo__sro_n1875;
wire CLOCK_slo__sro_n1922;


INV_X1 i_36 (.ZN (n_34), .A (Multiplier[30]));
INV_X2 i_35 (.ZN (n_33), .A (p_0[30]));
INV_X1 i_34 (.ZN (n_32), .A (n_30));
OAI33_X1 i_33 (.ZN (n_31), .A1 (n_32), .A2 (p_0[30]), .A3 (n_34), .B1 (n_30), .B2 (n_33), .B3 (Multiplier[30]));
XOR2_X1 i_32 (.Z (p_1[31]), .A (Multiplier[31]), .B (n_31));
OAI22_X1 i_31 (.ZN (n_0), .A1 (n_34), .A2 (p_0[30]), .B1 (Multiplier[30]), .B2 (n_33));
XNOR2_X1 i_0 (.ZN (p_1[30]), .A (n_0), .B (n_32));
XNOR2_X1 CLOCK_slo__sro_c1298 (.ZN (p_1[27]), .A (CLOCK_slo__sro_n1694), .B (n_27));
XNOR2_X2 slo__mro_c724 (.ZN (slo__mro_n875), .A (n_16), .B (Multiplier[16]));
OAI21_X1 CLOCK_slo__sro_c1404 (.ZN (CLOCK_slo__sro_n1809), .A (n_3), .B1 (p_0[3]), .B2 (Multiplier[3]));
INV_X1 slo__sro_c31 (.ZN (slo__sro_n88), .A (n_22));
FA_X1 i_26 (.CO (n_26), .S (p_1[25]), .A (Multiplier[25]), .B (p_0[25]), .CI (n_25));
FA_X1 i_25 (.CO (n_25), .S (p_1[24]), .A (Multiplier[24]), .B (p_0[24]), .CI (n_24));
NAND2_X1 slo__sro_c699 (.ZN (slo__sro_n848), .A1 (p_0[28]), .A2 (Multiplier[28]));
INV_X1 slo__sro_c45 (.ZN (slo__sro_n102), .A (n_11));
FA_X1 i_22 (.CO (n_22), .S (p_1[21]), .A (Multiplier[21]), .B (p_0[21]), .CI (n_21));
INV_X1 slo__sro_c217 (.ZN (slo__sro_n283), .A (p_0[1]));
INV_X1 slo__sro_c17 (.ZN (slo__sro_n75), .A (n_26));
NOR2_X1 slo__sro_c610 (.ZN (slo__sro_n751), .A1 (p_0[15]), .A2 (Multiplier[15]));
INV_X1 slo__sro_c181 (.ZN (slo__sro_n249), .A (p_0[12]));
NAND2_X1 slo__sro_c806 (.ZN (slo__sro_n993), .A1 (opt_ipoPP_0), .A2 (Multiplier[4]));
NAND2_X1 slo__sro_c687 (.ZN (slo__sro_n834), .A1 (p_0[23]), .A2 (Multiplier[23]));
FA_X1 i_15 (.CO (n_15), .S (p_1[14]), .A (Multiplier[14]), .B (p_0[14]), .CI (n_14));
FA_X1 i_14 (.CO (n_14), .S (p_1[13]), .A (Multiplier[13]), .B (p_0[13]), .CI (slo__sro_n246));
NAND2_X1 slo__sro_c195 (.ZN (slo__sro_n265), .A1 (p_0[20]), .A2 (Multiplier[20]));
INV_X1 slo__sro_c111 (.ZN (slo__sro_n171), .A (slo__sro_n991));
FA_X1 i_10 (.CO (n_10), .S (p_1[9]), .A (Multiplier[9]), .B (p_0[9]), .CI (n_9));
XNOR2_X1 CLOCK_slo__mro_c1122 (.ZN (CLOCK_slo__mro_n1455), .A (p_0[18]), .B (Multiplier[18]));
FA_X1 i_8 (.CO (n_8), .S (p_1[7]), .A (Multiplier[7]), .B (p_0[7]), .CI (n_7));
FA_X1 i_7 (.CO (n_7), .S (p_1[6]), .A (Multiplier[6]), .B (p_0[6]), .CI (slo__sro_n168));
INV_X1 slo__sro_c125 (.ZN (slo__sro_n188), .A (n_16));
INV_X1 CLOCK_slo__sro_c1084 (.ZN (CLOCK_slo__sro_n1422), .A (n_8));
NAND2_X1 CLOCK_slo__sro_c1467 (.ZN (CLOCK_slo__sro_n1874), .A1 (p_0[10]), .A2 (Multiplier[10]));
INV_X1 slo__L1_c1_c760 (.ZN (slo_n951), .A (p_0[17]));
NAND2_X1 slo__sro_c235 (.ZN (slo__sro_n299), .A1 (p_0[18]), .A2 (Multiplier[18]));
HA_X1 i_1 (.CO (n_1), .S (p_1[0]), .A (Multiplier[0]), .B (p_0[0]));
INV_X1 slo__sro_c3 (.ZN (slo__sro_n62), .A (n_19));
NAND2_X1 slo__sro_c4 (.ZN (slo__sro_n61), .A1 (p_0[19]), .A2 (Multiplier[19]));
NOR2_X1 slo__sro_c5 (.ZN (slo__sro_n60), .A1 (p_0[19]), .A2 (Multiplier[19]));
OAI21_X2 slo__sro_c6 (.ZN (n_20), .A (slo__sro_n61), .B1 (slo__sro_n62), .B2 (slo__sro_n60));
XNOR2_X2 slo__sro_c690 (.ZN (slo__sro_n832), .A (p_0[23]), .B (Multiplier[23]));
XNOR2_X2 slo__sro_c691 (.ZN (p_1[23]), .A (slo__sro_n832), .B (n_23));
NAND2_X1 slo__sro_c18 (.ZN (slo__sro_n74), .A1 (p_0[26]), .A2 (Multiplier[26]));
NOR2_X1 slo__sro_c19 (.ZN (slo__sro_n73), .A1 (p_0[26]), .A2 (Multiplier[26]));
OAI21_X1 slo__sro_c20 (.ZN (n_27), .A (slo__sro_n74), .B1 (slo__sro_n73), .B2 (slo__sro_n75));
INV_X2 slo__sro_c608 (.ZN (slo__sro_n753), .A (n_15));
NAND2_X1 slo__sro_c609 (.ZN (slo__sro_n752), .A1 (p_0[15]), .A2 (Multiplier[15]));
NAND2_X1 slo__sro_c32 (.ZN (slo__sro_n87), .A1 (p_0[22]), .A2 (Multiplier[22]));
OAI21_X2 slo__sro_c34 (.ZN (n_23), .A (slo__sro_n87), .B1 (slo__sro_n88), .B2 (CLOCK_slo__sro_n1922));
XNOR2_X2 slo__sro_c35 (.ZN (slo__sro_n85), .A (p_0[22]), .B (Multiplier[22]));
XNOR2_X2 slo__sro_c36 (.ZN (p_1[22]), .A (slo__sro_n85), .B (n_22));
NAND2_X1 slo__sro_c46 (.ZN (slo__sro_n101), .A1 (p_0[11]), .A2 (Multiplier[11]));
NOR2_X2 slo__sro_c47 (.ZN (slo__sro_n100), .A1 (p_0[11]), .A2 (Multiplier[11]));
OAI21_X2 slo__sro_c48 (.ZN (slo__sro_n99), .A (slo__sro_n101), .B1 (slo__sro_n102), .B2 (slo__sro_n100));
XNOR2_X1 slo__sro_c49 (.ZN (slo__sro_n98), .A (p_0[11]), .B (Multiplier[11]));
XNOR2_X1 slo__sro_c50 (.ZN (p_1[11]), .A (slo__sro_n98), .B (n_11));
NAND2_X1 slo__sro_c112 (.ZN (slo__sro_n170), .A1 (p_0[5]), .A2 (Multiplier[5]));
NOR2_X1 slo__sro_c113 (.ZN (slo__sro_n169), .A1 (p_0[5]), .A2 (Multiplier[5]));
OAI21_X1 slo__sro_c114 (.ZN (slo__sro_n168), .A (slo__sro_n170), .B1 (slo__sro_n171), .B2 (slo__sro_n169));
XNOR2_X2 slo__sro_c115 (.ZN (slo__sro_n167), .A (p_0[5]), .B (Multiplier[5]));
XNOR2_X2 slo__sro_c116 (.ZN (p_1[5]), .A (slo__sro_n167), .B (slo__sro_n991));
NAND2_X1 slo__sro_c126 (.ZN (slo__sro_n187), .A1 (p_0[16]), .A2 (Multiplier[16]));
NOR2_X1 CLOCK_slo__sro_c1086 (.ZN (CLOCK_slo__sro_n1420), .A1 (p_0[8]), .A2 (Multiplier[8]));
OAI21_X2 slo__sro_c128 (.ZN (slo__sro_n185), .A (slo__sro_n187), .B1 (slo__sro_n1234), .B2 (slo__sro_n188));
NAND2_X1 slo__sro_c732 (.ZN (slo__sro_n888), .A1 (p_0[2]), .A2 (Multiplier[2]));
OAI21_X1 slo__sro_c733 (.ZN (slo__sro_n887), .A (n_2), .B1 (p_0[2]), .B2 (Multiplier[2]));
NAND2_X1 slo__sro_c168 (.ZN (slo__sro_n231), .A1 (slo__sro_n185), .A2 (Multiplier[17]));
NOR2_X1 slo__sro_c169 (.ZN (slo__sro_n230), .A1 (slo__sro_n185), .A2 (Multiplier[17]));
OAI21_X1 slo__sro_c170 (.ZN (slo__sro_n229), .A (slo__sro_n231), .B1 (slo_n951), .B2 (slo__sro_n230));
XNOR2_X1 slo__sro_c171 (.ZN (slo__sro_n228), .A (slo__sro_n185), .B (Multiplier[17]));
XNOR2_X1 slo__sro_c172 (.ZN (p_1[17]), .A (slo__sro_n228), .B (p_0_17_PP_1));
NAND2_X1 slo__sro_c182 (.ZN (slo__sro_n248), .A1 (slo__sro_n99), .A2 (Multiplier[12]));
NOR2_X1 slo__sro_c183 (.ZN (slo__sro_n247), .A1 (slo__sro_n99), .A2 (Multiplier[12]));
OAI21_X1 slo__sro_c184 (.ZN (slo__sro_n246), .A (slo__sro_n248), .B1 (slo__sro_n247), .B2 (slo__sro_n249));
XNOR2_X1 slo__sro_c185 (.ZN (slo__sro_n245), .A (slo__sro_n99), .B (Multiplier[12]));
XNOR2_X1 slo__sro_c186 (.ZN (p_1[12]), .A (slo__sro_n245), .B (p_0[12]));
NAND2_X1 slo__sro_c689 (.ZN (n_24), .A1 (slo__sro_n834), .A2 (slo__sro_n833));
NAND2_X1 slo__sro_c197 (.ZN (slo__sro_n263), .A1 (n_20), .A2 (p_0[20]));
NAND3_X1 slo__sro_c198 (.ZN (n_21), .A1 (slo__sro_n263), .A2 (slo__mro_n826), .A3 (slo__sro_n265));
XNOR2_X2 slo__sro_c199 (.ZN (slo__sro_n262), .A (p_0[20]), .B (Multiplier[20]));
XNOR2_X1 slo__sro_c200 (.ZN (p_1[20]), .A (slo__sro_n262), .B (n_20));
NAND2_X1 slo__sro_c218 (.ZN (slo__sro_n282), .A1 (n_1), .A2 (Multiplier[1]));
NOR2_X1 slo__sro_c219 (.ZN (slo__sro_n281), .A1 (n_1), .A2 (Multiplier[1]));
OAI21_X1 slo__sro_c220 (.ZN (n_2), .A (slo__sro_n282), .B1 (slo__sro_n283), .B2 (slo__sro_n281));
XNOR2_X2 slo__sro_c221 (.ZN (slo__sro_n280), .A (n_1), .B (Multiplier[1]));
XNOR2_X1 slo__sro_c222 (.ZN (p_1[1]), .A (p_0[1]), .B (slo__sro_n280));
NAND2_X2 slo__sro_c237 (.ZN (n_19), .A1 (slo__sro_n299), .A2 (CLOCK_slo__sro_n1464));
OAI21_X1 CLOCK_slo__sro_c1130 (.ZN (CLOCK_slo__sro_n1464), .A (slo__sro_n229), .B1 (p_0[18]), .B2 (Multiplier[18]));
XNOR2_X1 CLOCK_slo__sro_c1203 (.ZN (p_1[26]), .A (slo__mro_n724), .B (n_26));
OAI21_X2 slo__sro_c611 (.ZN (n_16), .A (slo__sro_n752), .B1 (slo__sro_n753), .B2 (slo__sro_n751));
XNOR2_X1 slo__sro_c612 (.ZN (slo__sro_n750), .A (p_0[15]), .B (Multiplier[15]));
XNOR2_X1 slo__mro_c592 (.ZN (slo__mro_n724), .A (p_0[26]), .B (Multiplier[26]));
NAND2_X1 CLOCK_slo__sro_c1403 (.ZN (CLOCK_slo__sro_n1810), .A1 (p_0[3]), .A2 (Multiplier[3]));
XNOR2_X1 slo__sro_c613 (.ZN (p_1[15]), .A (slo__sro_n750), .B (n_15));
OAI21_X1 slo__sro_c688 (.ZN (slo__sro_n833), .A (n_23), .B1 (p_0[23]), .B2 (Multiplier[23]));
NAND2_X1 slo__mro_c683 (.ZN (slo__mro_n826), .A1 (n_20), .A2 (Multiplier[20]));
XNOR2_X2 slo__mro_c645 (.ZN (slo__mro_n796), .A (p_0[19]), .B (Multiplier[19]));
XNOR2_X2 slo__mro_c646 (.ZN (p_1[19]), .A (slo__mro_n796), .B (n_19));
OAI21_X1 slo__sro_c700 (.ZN (slo__sro_n847), .A (n_28), .B1 (p_0[28]), .B2 (Multiplier[28]));
NAND2_X1 slo__sro_c701 (.ZN (slo__sro_n846), .A1 (slo__sro_n847), .A2 (slo__sro_n848));
XNOR2_X2 slo__sro_c702 (.ZN (slo__sro_n845), .A (p_0[28]), .B (Multiplier[28]));
XNOR2_X2 slo__sro_c703 (.ZN (p_1[28]), .A (slo__sro_n845), .B (n_28));
XNOR2_X1 slo__mro_c725 (.ZN (p_1[16]), .A (slo__mro_n875), .B (p_0_16_PP_5));
NAND2_X1 slo__sro_c734 (.ZN (n_3), .A1 (slo__sro_n887), .A2 (slo__sro_n888));
XNOR2_X1 slo__sro_c735 (.ZN (slo__sro_n886), .A (p_0[2]), .B (Multiplier[2]));
XNOR2_X1 slo__sro_c736 (.ZN (p_1[2]), .A (slo__sro_n886), .B (n_2));
INV_X1 CLOCK_slo__sro_c1466 (.ZN (CLOCK_slo__sro_n1875), .A (n_10));
OAI21_X1 slo__sro_c807 (.ZN (slo__sro_n992), .A (CLOCK_slo__sro_n1808), .B1 (opt_ipoPP_0), .B2 (Multiplier[4]));
NAND2_X1 slo__sro_c808 (.ZN (slo__sro_n991), .A1 (slo__sro_n992), .A2 (slo__sro_n993));
XNOR2_X2 slo__sro_c809 (.ZN (slo__sro_n990), .A (p_0[4]), .B (Multiplier[4]));
XNOR2_X1 slo__sro_c810 (.ZN (p_1[4]), .A (slo__sro_n990), .B (CLOCK_slo__sro_n1808));
NAND2_X1 CLOCK_slo__sro_c1085 (.ZN (CLOCK_slo__sro_n1421), .A1 (p_0[8]), .A2 (Multiplier[8]));
NOR2_X2 slo__sro_c960 (.ZN (slo__sro_n1234), .A1 (p_0[16]), .A2 (Multiplier[16]));
OAI21_X2 CLOCK_slo__sro_c1087 (.ZN (n_9), .A (CLOCK_slo__sro_n1421), .B1 (CLOCK_slo__sro_n1422), .B2 (CLOCK_slo__sro_n1420));
XNOR2_X1 CLOCK_slo__sro_c1088 (.ZN (CLOCK_slo__sro_n1419), .A (p_0[8]), .B (Multiplier[8]));
XNOR2_X1 CLOCK_slo__sro_c1089 (.ZN (p_1[8]), .A (CLOCK_slo__sro_n1419), .B (n_8));
XNOR2_X1 CLOCK_slo__mro_c1123 (.ZN (p_1[18]), .A (CLOCK_slo__mro_n1455), .B (slo__sro_n229));
NAND2_X1 CLOCK_slo__sro_c1294 (.ZN (CLOCK_slo__sro_n1696), .A1 (p_0[27]), .A2 (Multiplier[27]));
OAI21_X1 CLOCK_slo__sro_c1295 (.ZN (CLOCK_slo__sro_n1695), .A (n_27), .B1 (p_0[27]), .B2 (Multiplier[27]));
NAND2_X1 CLOCK_slo__sro_c1296 (.ZN (n_28), .A1 (CLOCK_slo__sro_n1695), .A2 (CLOCK_slo__sro_n1696));
XNOR2_X1 CLOCK_slo__sro_c1297 (.ZN (CLOCK_slo__sro_n1694), .A (p_0[27]), .B (Multiplier[27]));
INV_X1 CLOCK_slo__sro_c1151 (.ZN (CLOCK_slo__sro_n1489), .A (slo__sro_n846));
NAND2_X1 CLOCK_slo__sro_c1152 (.ZN (CLOCK_slo__sro_n1488), .A1 (p_0[29]), .A2 (Multiplier[29]));
NOR2_X1 CLOCK_slo__sro_c1153 (.ZN (CLOCK_slo__sro_n1487), .A1 (p_0[29]), .A2 (Multiplier[29]));
OAI21_X1 CLOCK_slo__sro_c1154 (.ZN (n_30), .A (CLOCK_slo__sro_n1488), .B1 (CLOCK_slo__sro_n1489), .B2 (CLOCK_slo__sro_n1487));
XNOR2_X1 CLOCK_slo__sro_c1155 (.ZN (CLOCK_slo__sro_n1486), .A (p_0[29]), .B (Multiplier[29]));
XNOR2_X1 CLOCK_slo__sro_c1156 (.ZN (p_1[29]), .A (CLOCK_slo__sro_n1486), .B (slo__sro_n846));
NAND2_X1 CLOCK_slo__sro_c1405 (.ZN (CLOCK_slo__sro_n1808), .A1 (CLOCK_slo__sro_n1810), .A2 (CLOCK_slo__sro_n1809));
XNOR2_X1 CLOCK_slo__sro_c1406 (.ZN (CLOCK_slo__sro_n1807), .A (p_0[3]), .B (Multiplier[3]));
XNOR2_X1 CLOCK_slo__sro_c1407 (.ZN (p_1[3]), .A (CLOCK_slo__sro_n1807), .B (n_3));
NOR2_X1 CLOCK_slo__sro_c1468 (.ZN (CLOCK_slo__sro_n1873), .A1 (p_0[10]), .A2 (Multiplier[10]));
OAI21_X2 CLOCK_slo__sro_c1469 (.ZN (n_11), .A (CLOCK_slo__sro_n1874), .B1 (CLOCK_slo__sro_n1873), .B2 (CLOCK_slo__sro_n1875));
XNOR2_X2 CLOCK_slo__sro_c1470 (.ZN (CLOCK_slo__sro_n1872), .A (p_0[10]), .B (Multiplier[10]));
XNOR2_X2 CLOCK_slo__sro_c1471 (.ZN (p_1[10]), .A (CLOCK_slo__sro_n1872), .B (n_10));
NOR2_X2 CLOCK_slo__sro_c1514 (.ZN (CLOCK_slo__sro_n1922), .A1 (p_0[22]), .A2 (Multiplier[22]));

endmodule //datapath__0_201

module datapath__0_197 (opt_ipoPP_1, p_0, p_1, p_2);

output [31:0] p_2;
input [31:0] p_0;
input [31:0] p_1;
input opt_ipoPP_1;
wire slo__sro_n1043;
wire slo__sro_n1010;
wire n_1;
wire n_2;
wire n_3;
wire n_4;
wire n_5;
wire n_6;
wire n_7;
wire n_8;
wire n_9;
wire n_10;
wire n_11;
wire n_12;
wire n_13;
wire n_14;
wire n_15;
wire n_16;
wire slo__sro_n1011;
wire n_18;
wire n_19;
wire n_20;
wire n_21;
wire n_22;
wire n_23;
wire n_24;
wire n_25;
wire n_26;
wire n_27;
wire n_30;
wire n_32;
wire n_0;
wire n_34;
wire n_33;
wire slo__sro_n272;
wire slo__sro_n273;
wire slo__sro_n274;
wire slo__sro_n275;
wire slo__sro_n259;
wire slo__sro_n260;
wire slo__sro_n261;
wire slo__sro_n262;
wire slo__sro_n300;
wire slo__sro_n301;
wire slo__sro_n302;
wire slo__sro_n303;
wire slo__sro_n743;
wire slo__sro_n744;
wire slo__sro_n745;
wire slo__sro_n746;
wire slo__sro_n578;
wire slo__sro_n579;
wire slo__sro_n580;
wire slo__sro_n581;
wire slo__sro_n582;
wire slo__sro_n1012;
wire slo__sro_n1013;
wire slo__sro_n1044;
wire slo__sro_n1045;
wire slo__sro_n144;
wire slo__sro_n145;
wire slo__sro_n146;
wire slo__sro_n147;
wire slo__sro_n1046;
wire slo__sro_n1047;
wire slo__sro_n1057;
wire slo__sro_n1058;
wire slo__sro_n375;
wire slo__sro_n376;
wire slo__sro_n377;
wire slo__sro_n378;
wire slo__sro_n1059;
wire slo__sro_n1060;
wire slo__sro_n1061;
wire CLOCK_slo__sro_n1292;
wire CLOCK_slo__sro_n1293;
wire CLOCK_slo__sro_n1294;
wire CLOCK_slo__sro_n1295;
wire slo__sro_n1114;
wire slo__sro_n1115;
wire slo__sro_n1116;
wire slo__sro_n1117;
wire CLOCK_slo__sro_n1373;
wire CLOCK_slo__sro_n1374;
wire CLOCK_slo__sro_n1375;
wire CLOCK_slo__sro_n1376;
wire CLOCK_slo__sro_n1461;
wire CLOCK_slo__sro_n1462;
wire CLOCK_slo__sro_n1463;
wire CLOCK_slo__sro_n1464;
wire CLOCK_slo__sro_n1699;
wire CLOCK_slo__sro_n1700;
wire CLOCK_slo__sro_n1701;
wire CLOCK_slo__sro_n1702;
wire CLOCK_slo__sro_n1703;
wire CLOCK_slo__sro_n1663;
wire CLOCK_slo__sro_n1664;
wire CLOCK_slo__sro_n1665;
wire CLOCK_slo__sro_n1666;


INV_X1 i_36 (.ZN (n_34), .A (p_0[30]));
INV_X1 i_35 (.ZN (n_33), .A (p_1[30]));
INV_X2 i_34 (.ZN (n_32), .A (n_30));
INV_X1 slo__sro_c805 (.ZN (slo__sro_n1061), .A (CLOCK_slo__sro_n1700));
XOR2_X1 i_32 (.Z (p_2[31]), .A (p_0[31]), .B (slo__sro_n1043));
OAI22_X1 i_31 (.ZN (n_0), .A1 (n_34), .A2 (p_1[30]), .B1 (p_0[30]), .B2 (n_33));
XNOR2_X1 i_0 (.ZN (p_2[30]), .A (n_32), .B (n_0));
FA_X1 i_30 (.CO (n_30), .S (p_2[29]), .A (p_0[29]), .B (p_1[29]), .CI (slo__sro_n1058));
INV_X1 CLOCK_slo__sro_c938 (.ZN (CLOCK_slo__sro_n1295), .A (n_4));
FA_X1 i_27 (.CO (n_27), .S (p_2[26]), .A (p_0[26]), .B (p_1[26]), .CI (n_26));
FA_X1 i_26 (.CO (n_26), .S (p_2[25]), .A (p_0[25]), .B (p_1[25]), .CI (n_25));
FA_X1 i_25 (.CO (n_25), .S (p_2[24]), .A (p_0[24]), .B (p_1[24]), .CI (n_24));
NAND2_X1 CLOCK_slo__sro_c1026 (.ZN (CLOCK_slo__sro_n1375), .A1 (p_1[15]), .A2 (p_0[15]));
INV_X1 slo__sro_c793 (.ZN (slo__sro_n1047), .A (n_34));
FA_X1 i_22 (.CO (n_22), .S (p_2[21]), .A (p_0[21]), .B (p_1[21]), .CI (n_21));
INV_X1 slo__sro_c233 (.ZN (slo__sro_n303), .A (p_1[1]));
FA_X1 i_20 (.CO (n_20), .S (p_2[19]), .A (p_0[19]), .B (p_1[19]), .CI (n_19));
FA_X1 i_19 (.CO (n_19), .S (p_2[18]), .A (p_0[18]), .B (p_1[18]), .CI (n_18));
INV_X1 CLOCK_slo__sro_c1301 (.ZN (CLOCK_slo__sro_n1703), .A (n_27));
XNOR2_X1 slo__sro_c578 (.ZN (p_2[7]), .A (slo__sro_n743), .B (n_7));
NAND2_X1 slo__sro_c234 (.ZN (slo__sro_n302), .A1 (n_1), .A2 (p_0[1]));
FA_X1 i_14 (.CO (n_14), .S (p_2[13]), .A (p_0[13]), .B (p_1[13]), .CI (n_13));
XNOR2_X1 slo__sro_c810 (.ZN (p_2[28]), .A (slo__sro_n1057), .B (CLOCK_slo__sro_n1700));
NOR2_X4 slo__sro_c807 (.ZN (slo__sro_n1059), .A1 (opt_ipoPP_1), .A2 (p_0[28]));
FA_X1 i_10 (.CO (n_10), .S (p_2[9]), .A (p_0[9]), .B (p_1[9]), .CI (n_9));
FA_X1 i_9 (.CO (n_9), .S (p_2[8]), .A (p_0[8]), .B (p_1[8]), .CI (n_8));
NAND2_X1 slo__sro_c765 (.ZN (slo__sro_n1012), .A1 (p_1[22]), .A2 (p_0[22]));
FA_X1 i_7 (.CO (n_7), .S (p_2[6]), .A (p_0[6]), .B (p_1[6]), .CI (n_6));
FA_X1 i_6 (.CO (n_6), .S (p_2[5]), .A (p_0[5]), .B (p_1[5]), .CI (n_5));
INV_X1 CLOCK_slo__sro_c1025 (.ZN (CLOCK_slo__sro_n1376), .A (n_15));
FA_X1 i_4 (.CO (n_4), .S (p_2[3]), .A (p_0[3]), .B (p_1[3]), .CI (n_3));
FA_X1 i_3 (.CO (n_3), .S (p_2[2]), .A (p_0[2]), .B (p_1[2]), .CI (n_2));
INV_X1 slo__sro_c764 (.ZN (slo__sro_n1013), .A (n_22));
HA_X1 i_1 (.CO (n_1), .S (p_2[0]), .A (p_0[0]), .B (p_1[0]));
INV_X1 slo__sro_c204 (.ZN (slo__sro_n275), .A (n_20));
NAND2_X1 slo__sro_c205 (.ZN (slo__sro_n274), .A1 (p_1[20]), .A2 (p_0[20]));
NOR2_X1 slo__sro_c206 (.ZN (slo__sro_n273), .A1 (p_1[20]), .A2 (p_0[20]));
OAI21_X1 slo__sro_c207 (.ZN (n_21), .A (slo__sro_n274), .B1 (slo__sro_n275), .B2 (slo__sro_n273));
XNOR2_X1 slo__sro_c208 (.ZN (slo__sro_n272), .A (p_1[20]), .B (p_0[20]));
XNOR2_X1 slo__sro_c209 (.ZN (p_2[20]), .A (n_20), .B (slo__sro_n272));
INV_X1 slo__sro_c190 (.ZN (slo__sro_n262), .A (n_14));
NAND2_X1 slo__sro_c191 (.ZN (slo__sro_n261), .A1 (p_1[14]), .A2 (p_0[14]));
NOR2_X1 slo__sro_c192 (.ZN (slo__sro_n260), .A1 (p_1[14]), .A2 (p_0[14]));
OAI21_X1 slo__sro_c193 (.ZN (n_15), .A (slo__sro_n261), .B1 (slo__sro_n262), .B2 (slo__sro_n260));
XNOR2_X1 slo__sro_c194 (.ZN (slo__sro_n259), .A (p_1[14]), .B (p_0[14]));
XNOR2_X1 slo__sro_c195 (.ZN (p_2[14]), .A (slo__sro_n259), .B (n_14));
NOR2_X1 slo__sro_c235 (.ZN (slo__sro_n301), .A1 (n_1), .A2 (p_0[1]));
OAI21_X1 slo__sro_c236 (.ZN (n_2), .A (slo__sro_n302), .B1 (slo__sro_n303), .B2 (slo__sro_n301));
XNOR2_X1 slo__sro_c237 (.ZN (slo__sro_n300), .A (n_1), .B (p_0[1]));
XNOR2_X1 slo__sro_c238 (.ZN (p_2[1]), .A (p_1[1]), .B (slo__sro_n300));
INV_X1 slo__sro_c573 (.ZN (slo__sro_n746), .A (n_7));
NAND2_X1 slo__sro_c574 (.ZN (slo__sro_n745), .A1 (p_1[7]), .A2 (p_0[7]));
NOR2_X1 slo__sro_c575 (.ZN (slo__sro_n744), .A1 (p_1[7]), .A2 (p_0[7]));
OAI21_X1 slo__sro_c576 (.ZN (n_8), .A (slo__sro_n745), .B1 (slo__sro_n746), .B2 (slo__sro_n744));
XNOR2_X1 slo__sro_c577 (.ZN (slo__sro_n743), .A (p_1[7]), .B (p_0[7]));
INV_X1 slo__sro_c459 (.ZN (slo__sro_n582), .A (n_16));
NAND2_X1 slo__sro_c460 (.ZN (slo__sro_n581), .A1 (p_0[16]), .A2 (p_1[16]));
NOR2_X1 slo__sro_c461 (.ZN (slo__sro_n580), .A1 (p_1[16]), .A2 (p_0[16]));
OAI21_X2 slo__sro_c462 (.ZN (slo__sro_n579), .A (slo__sro_n581), .B1 (slo__sro_n582), .B2 (slo__sro_n580));
XNOR2_X1 slo__sro_c463 (.ZN (slo__sro_n578), .A (p_1[16]), .B (p_0[16]));
XNOR2_X1 slo__sro_c464 (.ZN (p_2[16]), .A (slo__sro_n578), .B (n_16));
NOR2_X1 slo__sro_c766 (.ZN (slo__sro_n1011), .A1 (p_1[22]), .A2 (p_0[22]));
OAI21_X1 slo__sro_c767 (.ZN (n_23), .A (slo__sro_n1012), .B1 (slo__sro_n1013), .B2 (slo__sro_n1011));
XNOR2_X1 slo__sro_c768 (.ZN (slo__sro_n1010), .A (p_1[22]), .B (p_0[22]));
XNOR2_X1 slo__sro_c769 (.ZN (p_2[22]), .A (slo__sro_n1010), .B (n_22));
INV_X1 slo__sro_c794 (.ZN (slo__sro_n1046), .A (p_1[30]));
OR2_X1 slo__sro_c795 (.ZN (slo__sro_n1045), .A1 (n_33), .A2 (p_0[30]));
NAND2_X1 slo__sro_c796 (.ZN (slo__sro_n1044), .A1 (slo__sro_n1046), .A2 (slo__sro_n1047));
OAI22_X1 slo__sro_c797 (.ZN (slo__sro_n1043), .A1 (n_32), .A2 (slo__sro_n1044), .B1 (n_30), .B2 (slo__sro_n1045));
NAND2_X1 slo__sro_c806 (.ZN (slo__sro_n1060), .A1 (opt_ipoPP_1), .A2 (p_0[28]));
INV_X1 slo__sro_c85 (.ZN (slo__sro_n147), .A (n_11));
NAND2_X1 slo__sro_c86 (.ZN (slo__sro_n146), .A1 (p_1[11]), .A2 (p_0[11]));
NOR2_X1 slo__sro_c87 (.ZN (slo__sro_n145), .A1 (p_1[11]), .A2 (p_0[11]));
OAI21_X1 slo__sro_c88 (.ZN (n_12), .A (slo__sro_n146), .B1 (slo__sro_n147), .B2 (slo__sro_n145));
XNOR2_X1 slo__sro_c89 (.ZN (slo__sro_n144), .A (p_1[11]), .B (p_0[11]));
XNOR2_X1 slo__sro_c90 (.ZN (p_2[11]), .A (slo__sro_n144), .B (n_11));
OAI21_X1 slo__sro_c808 (.ZN (slo__sro_n1058), .A (slo__sro_n1060), .B1 (slo__sro_n1059), .B2 (slo__sro_n1061));
XNOR2_X1 slo__sro_c809 (.ZN (slo__sro_n1057), .A (p_1[28]), .B (p_0[28]));
INV_X1 slo__sro_c314 (.ZN (slo__sro_n378), .A (n_12));
NAND2_X1 slo__sro_c315 (.ZN (slo__sro_n377), .A1 (p_1[12]), .A2 (p_0[12]));
NOR2_X1 slo__sro_c316 (.ZN (slo__sro_n376), .A1 (p_1[12]), .A2 (p_0[12]));
OAI21_X1 slo__sro_c317 (.ZN (n_13), .A (slo__sro_n377), .B1 (slo__sro_n378), .B2 (slo__sro_n376));
XNOR2_X1 slo__sro_c318 (.ZN (slo__sro_n375), .A (p_1[12]), .B (p_0[12]));
XNOR2_X1 slo__sro_c319 (.ZN (p_2[12]), .A (slo__sro_n375), .B (n_12));
NAND2_X1 CLOCK_slo__sro_c939 (.ZN (CLOCK_slo__sro_n1294), .A1 (p_0[4]), .A2 (p_1[4]));
NOR2_X1 CLOCK_slo__sro_c940 (.ZN (CLOCK_slo__sro_n1293), .A1 (p_1[4]), .A2 (p_0[4]));
OAI21_X1 CLOCK_slo__sro_c941 (.ZN (n_5), .A (CLOCK_slo__sro_n1294), .B1 (CLOCK_slo__sro_n1295), .B2 (CLOCK_slo__sro_n1293));
XNOR2_X1 CLOCK_slo__sro_c942 (.ZN (CLOCK_slo__sro_n1292), .A (p_1[4]), .B (p_0[4]));
XNOR2_X1 CLOCK_slo__sro_c943 (.ZN (p_2[4]), .A (CLOCK_slo__sro_n1292), .B (n_4));
INV_X1 slo__sro_c849 (.ZN (slo__sro_n1117), .A (n_23));
NAND2_X1 slo__sro_c850 (.ZN (slo__sro_n1116), .A1 (p_1[23]), .A2 (p_0[23]));
NOR2_X1 slo__sro_c851 (.ZN (slo__sro_n1115), .A1 (p_1[23]), .A2 (p_0[23]));
OAI21_X1 slo__sro_c852 (.ZN (n_24), .A (slo__sro_n1116), .B1 (slo__sro_n1117), .B2 (slo__sro_n1115));
XNOR2_X1 slo__sro_c853 (.ZN (slo__sro_n1114), .A (p_1[23]), .B (p_0[23]));
XNOR2_X1 slo__sro_c854 (.ZN (p_2[23]), .A (slo__sro_n1114), .B (n_23));
NOR2_X1 CLOCK_slo__sro_c1027 (.ZN (CLOCK_slo__sro_n1374), .A1 (p_1[15]), .A2 (p_0[15]));
OAI21_X1 CLOCK_slo__sro_c1028 (.ZN (n_16), .A (CLOCK_slo__sro_n1375), .B1 (CLOCK_slo__sro_n1376), .B2 (CLOCK_slo__sro_n1374));
XNOR2_X1 CLOCK_slo__sro_c1029 (.ZN (CLOCK_slo__sro_n1373), .A (p_1[15]), .B (p_0[15]));
XNOR2_X2 CLOCK_slo__sro_c1030 (.ZN (p_2[15]), .A (CLOCK_slo__sro_n1373), .B (n_15));
NAND2_X1 CLOCK_slo__sro_c1106 (.ZN (CLOCK_slo__sro_n1464), .A1 (p_1[17]), .A2 (p_0[17]));
NAND2_X1 CLOCK_slo__sro_c1107 (.ZN (CLOCK_slo__sro_n1463), .A1 (slo__sro_n579), .A2 (p_0[17]));
NAND2_X1 CLOCK_slo__sro_c1108 (.ZN (CLOCK_slo__sro_n1462), .A1 (p_1[17]), .A2 (slo__sro_n579));
NAND3_X1 CLOCK_slo__sro_c1109 (.ZN (n_18), .A1 (CLOCK_slo__sro_n1462), .A2 (CLOCK_slo__sro_n1464), .A3 (CLOCK_slo__sro_n1463));
XNOR2_X1 CLOCK_slo__sro_c1110 (.ZN (CLOCK_slo__sro_n1461), .A (slo__sro_n579), .B (p_0[17]));
XNOR2_X1 CLOCK_slo__sro_c1111 (.ZN (p_2[17]), .A (CLOCK_slo__sro_n1461), .B (p_1[17]));
NAND2_X1 CLOCK_slo__sro_c1302 (.ZN (CLOCK_slo__sro_n1702), .A1 (p_0[27]), .A2 (p_1[27]));
NOR2_X1 CLOCK_slo__sro_c1303 (.ZN (CLOCK_slo__sro_n1701), .A1 (p_1[27]), .A2 (p_0[27]));
OAI21_X1 CLOCK_slo__sro_c1304 (.ZN (CLOCK_slo__sro_n1700), .A (CLOCK_slo__sro_n1702)
    , .B1 (CLOCK_slo__sro_n1703), .B2 (CLOCK_slo__sro_n1701));
XNOR2_X1 CLOCK_slo__sro_c1305 (.ZN (CLOCK_slo__sro_n1699), .A (p_1[27]), .B (p_0[27]));
XNOR2_X1 CLOCK_slo__sro_c1306 (.ZN (p_2[27]), .A (CLOCK_slo__sro_n1699), .B (n_27));
INV_X1 CLOCK_slo__sro_c1268 (.ZN (CLOCK_slo__sro_n1666), .A (n_10));
NAND2_X1 CLOCK_slo__sro_c1269 (.ZN (CLOCK_slo__sro_n1665), .A1 (p_0[10]), .A2 (p_1[10]));
NOR2_X1 CLOCK_slo__sro_c1270 (.ZN (CLOCK_slo__sro_n1664), .A1 (p_1[10]), .A2 (p_0[10]));
OAI21_X1 CLOCK_slo__sro_c1271 (.ZN (n_11), .A (CLOCK_slo__sro_n1665), .B1 (CLOCK_slo__sro_n1666), .B2 (CLOCK_slo__sro_n1664));
XNOR2_X1 CLOCK_slo__sro_c1272 (.ZN (CLOCK_slo__sro_n1663), .A (p_1[10]), .B (p_0[10]));
XNOR2_X1 CLOCK_slo__sro_c1273 (.ZN (p_2[10]), .A (n_10), .B (CLOCK_slo__sro_n1663));

endmodule //datapath__0_197

module datapath__0_196 (opt_ipoPP_1, Multiplier, p_0, p_1);

output [31:0] p_1;
input [31:0] Multiplier;
input [31:0] p_0;
input opt_ipoPP_1;
wire slo__sro_n464;
wire slo__mro_n851;
wire CLOCK_slo__sro_n1760;
wire n_1;
wire n_2;
wire n_3;
wire n_5;
wire n_6;
wire n_7;
wire n_8;
wire n_9;
wire n_10;
wire n_11;
wire n_12;
wire n_13;
wire n_14;
wire n_16;
wire n_18;
wire n_19;
wire n_21;
wire slo__sro_n880;
wire n_23;
wire n_25;
wire n_27;
wire n_28;
wire n_30;
wire n_32;
wire n_0;
wire n_34;
wire n_33;
wire n_31;
wire slo__sro_n57;
wire slo__sro_n58;
wire slo__sro_n59;
wire slo__sro_n60;
wire slo__sro_n61;
wire slo__sro_n74;
wire slo__sro_n75;
wire slo__sro_n76;
wire slo__sro_n77;
wire slo__sro_n87;
wire slo__sro_n88;
wire slo__sro_n89;
wire slo__sro_n90;
wire slo__sro_n91;
wire slo__sro_n159;
wire slo__sro_n160;
wire slo__sro_n161;
wire slo__sro_n162;
wire slo__sro_n163;
wire CLOCK_slo__sro_n1759;
wire slo__sro_n132;
wire slo__sro_n133;
wire slo__sro_n134;
wire slo__sro_n176;
wire slo__sro_n177;
wire slo__sro_n178;
wire slo__sro_n179;
wire slo__sro_n180;
wire slo__sro_n194;
wire slo__sro_n195;
wire slo__sro_n196;
wire slo__sro_n197;
wire slo__sro_n210;
wire slo__sro_n211;
wire slo__sro_n212;
wire slo__sro_n213;
wire slo__sro_n223;
wire slo__sro_n224;
wire slo__sro_n225;
wire slo__sro_n226;
wire slo__sro_n238;
wire slo__sro_n239;
wire slo__sro_n240;
wire slo__sro_n241;
wire slo__sro_n242;
wire slo__sro_n277;
wire slo__sro_n278;
wire slo__sro_n279;
wire slo__sro_n280;
wire slo__sro_n281;
wire slo__sro_n461;
wire slo__sro_n462;
wire slo__sro_n463;
wire slo__sro_n306;
wire slo__sro_n307;
wire slo__sro_n308;
wire slo__sro_n309;
wire slo__sro_n559;
wire slo__sro_n560;
wire slo__sro_n561;
wire slo__sro_n562;
wire slo__sro_n646;
wire slo__sro_n647;
wire slo__sro_n648;
wire slo__sro_n649;
wire slo__sro_n650;
wire slo__sro_n881;
wire slo__sro_n882;
wire slo__sro_n908;
wire slo__sro_n909;
wire slo__sro_n910;
wire slo__sro_n911;
wire CLOCK_slo__mro_n1383;
wire CLOCK_slo__sro_n1335;
wire CLOCK_slo__sro_n1336;
wire CLOCK_slo__sro_n1337;
wire CLOCK_slo__sro_n1523;
wire CLOCK_slo__sro_n1524;
wire CLOCK_slo__sro_n1525;
wire CLOCK_slo__sro_n1526;


INV_X1 i_36 (.ZN (n_34), .A (Multiplier[30]));
INV_X1 i_35 (.ZN (n_33), .A (p_0[30]));
INV_X1 i_34 (.ZN (n_32), .A (n_30));
XOR2_X1 i_32 (.Z (p_1[31]), .A (Multiplier[31]), .B (n_31));
OAI22_X1 i_31 (.ZN (n_0), .A1 (n_34), .A2 (p_0[30]), .B1 (Multiplier[30]), .B2 (n_33));
XNOR2_X1 i_0 (.ZN (p_1[30]), .A (n_32), .B (n_0));
FA_X1 i_30 (.CO (n_30), .S (p_1[29]), .A (Multiplier[29]), .B (p_0[29]), .CI (slo__sro_n194));
INV_X1 slo__sro_c138 (.ZN (slo__sro_n213), .A (p_0[1]));
INV_X1 slo__sro_c463 (.ZN (slo__sro_n650), .A (n_16));
FA_X1 i_27 (.CO (n_27), .S (p_1[26]), .A (Multiplier[26]), .B (p_0[26]), .CI (slo__sro_n278));
NAND2_X1 slo__sro_c402 (.ZN (slo__sro_n561), .A1 (p_0[27]), .A2 (Multiplier[27]));
FA_X1 i_25 (.CO (n_25), .S (p_1[24]), .A (Multiplier[24]), .B (p_0[24]), .CI (slo__sro_n58));
INV_X1 slo__sro_c15 (.ZN (slo__sro_n77), .A (n_11));
INV_X1 slo__sro_c626 (.ZN (slo__sro_n911), .A (n_9));
INV_X1 slo__sro_c124 (.ZN (slo__sro_n197), .A (n_28));
OAI22_X1 CLOCK_slo__sro_c1215 (.ZN (n_31), .A1 (n_32), .A2 (CLOCK_slo__sro_n1759)
    , .B1 (CLOCK_slo__sro_n1760), .B2 (n_30));
INV_X1 slo__sro_c96 (.ZN (slo__sro_n163), .A (n_14));
FA_X1 i_19 (.CO (n_19), .S (p_1[18]), .A (Multiplier[18]), .B (p_0[18]), .CI (n_18));
XNOR2_X1 slo__sro_c334 (.ZN (p_1[10]), .A (slo__sro_n461), .B (n_10));
XNOR2_X1 slo__mro_c585 (.ZN (p_1[28]), .A (slo__mro_n851), .B (p_0[28]));
FA_X1 i_16 (.CO (n_16), .S (p_1[15]), .A (Multiplier[15]), .B (p_0[15]), .CI (slo__sro_n160));
INV_X1 slo__sro_c110 (.ZN (slo__sro_n180), .A (n_21));
FA_X1 i_14 (.CO (n_14), .S (p_1[13]), .A (Multiplier[13]), .B (p_0[13]), .CI (n_13));
FA_X1 i_13 (.CO (n_13), .S (p_1[12]), .A (Multiplier[12]), .B (p_0[12]), .CI (n_12));
INV_X1 slo__sro_c29 (.ZN (slo__sro_n91), .A (n_19));
XNOR2_X2 slo__mro_c584 (.ZN (slo__mro_n851), .A (n_28), .B (Multiplier[28]));
INV_X1 CLOCK_slo__sro_c1009 (.ZN (CLOCK_slo__sro_n1526), .A (slo__sro_n88));
FA_X1 i_9 (.CO (n_9), .S (p_1[8]), .A (Multiplier[8]), .B (p_0[8]), .CI (n_8));
INV_X1 slo__sro_c166 (.ZN (slo__sro_n242), .A (n_3));
NAND2_X1 slo__sro_c111 (.ZN (slo__sro_n179), .A1 (p_0[21]), .A2 (Multiplier[21]));
XNOR2_X2 CLOCK_slo__mro_c896 (.ZN (CLOCK_slo__mro_n1383), .A (n_6), .B (Multiplier[6]));
FA_X1 i_5 (.CO (n_5), .S (p_1[4]), .A (Multiplier[4]), .B (p_0[4]), .CI (slo__sro_n239));
INV_X1 slo__sro_c200 (.ZN (slo__sro_n281), .A (n_25));
FA_X1 i_3 (.CO (n_3), .S (p_1[2]), .A (Multiplier[2]), .B (p_0[2]), .CI (n_2));
INV_X1 slo__sro_c152 (.ZN (slo__sro_n226), .A (p_0[7]));
HA_X1 i_1 (.CO (n_1), .S (p_1[0]), .A (Multiplier[0]), .B (p_0[0]));
INV_X1 slo__sro_c1 (.ZN (slo__sro_n61), .A (n_23));
NAND2_X1 slo__sro_c2 (.ZN (slo__sro_n60), .A1 (p_0[23]), .A2 (Multiplier[23]));
NOR2_X1 slo__sro_c3 (.ZN (slo__sro_n59), .A1 (p_0[23]), .A2 (Multiplier[23]));
OAI21_X1 slo__sro_c4 (.ZN (slo__sro_n58), .A (slo__sro_n60), .B1 (slo__sro_n59), .B2 (slo__sro_n61));
XNOR2_X2 slo__sro_c5 (.ZN (slo__sro_n57), .A (p_0[23]), .B (Multiplier[23]));
XNOR2_X2 slo__sro_c6 (.ZN (p_1[23]), .A (slo__sro_n57), .B (n_23));
NAND2_X1 slo__sro_c16 (.ZN (slo__sro_n76), .A1 (p_0[11]), .A2 (Multiplier[11]));
NOR2_X1 slo__sro_c17 (.ZN (slo__sro_n75), .A1 (p_0[11]), .A2 (Multiplier[11]));
OAI21_X1 slo__sro_c18 (.ZN (n_12), .A (slo__sro_n76), .B1 (slo__sro_n77), .B2 (slo__sro_n75));
XNOR2_X1 slo__sro_c19 (.ZN (slo__sro_n74), .A (p_0[11]), .B (Multiplier[11]));
XNOR2_X1 slo__sro_c20 (.ZN (p_1[11]), .A (slo__sro_n74), .B (n_11));
NAND2_X1 slo__sro_c30 (.ZN (slo__sro_n90), .A1 (p_0[19]), .A2 (Multiplier[19]));
NOR2_X1 slo__sro_c31 (.ZN (slo__sro_n89), .A1 (p_0[19]), .A2 (Multiplier[19]));
OAI21_X1 slo__sro_c32 (.ZN (slo__sro_n88), .A (slo__sro_n90), .B1 (slo__sro_n91), .B2 (slo__sro_n89));
XNOR2_X1 slo__sro_c33 (.ZN (slo__sro_n87), .A (p_0[19]), .B (Multiplier[19]));
XNOR2_X1 slo__sro_c34 (.ZN (p_1[19]), .A (slo__sro_n87), .B (n_19));
NAND2_X1 slo__sro_c97 (.ZN (slo__sro_n162), .A1 (p_0[14]), .A2 (Multiplier[14]));
NOR2_X1 slo__sro_c98 (.ZN (slo__sro_n161), .A1 (p_0[14]), .A2 (Multiplier[14]));
OAI21_X1 slo__sro_c99 (.ZN (slo__sro_n160), .A (slo__sro_n162), .B1 (slo__sro_n163), .B2 (slo__sro_n161));
XNOR2_X1 slo__sro_c100 (.ZN (slo__sro_n159), .A (p_0[14]), .B (Multiplier[14]));
XNOR2_X1 slo__sro_c101 (.ZN (p_1[14]), .A (slo__sro_n159), .B (n_14));
INV_X1 slo__sro_c69 (.ZN (slo__sro_n134), .A (n_6));
NAND2_X1 slo__sro_c70 (.ZN (slo__sro_n133), .A1 (p_0[6]), .A2 (Multiplier[6]));
NOR2_X1 slo__sro_c71 (.ZN (slo__sro_n132), .A1 (p_0[6]), .A2 (Multiplier[6]));
OAI21_X2 slo__sro_c72 (.ZN (n_7), .A (slo__sro_n133), .B1 (slo__sro_n132), .B2 (slo__sro_n134));
OR2_X1 CLOCK_slo__sro_c1213 (.ZN (CLOCK_slo__sro_n1760), .A1 (n_33), .A2 (Multiplier[30]));
XNOR2_X1 CLOCK_slo__sro_c972 (.ZN (p_1[3]), .A (slo__sro_n238), .B (n_3));
NOR2_X1 slo__sro_c112 (.ZN (slo__sro_n178), .A1 (p_0[21]), .A2 (Multiplier[21]));
OAI21_X1 slo__sro_c113 (.ZN (slo__sro_n177), .A (slo__sro_n179), .B1 (slo__sro_n178), .B2 (slo__sro_n180));
XNOR2_X1 slo__sro_c114 (.ZN (slo__sro_n176), .A (p_0[21]), .B (Multiplier[21]));
XNOR2_X1 slo__sro_c115 (.ZN (p_1[21]), .A (slo__sro_n176), .B (n_21));
NAND2_X1 slo__sro_c125 (.ZN (slo__sro_n196), .A1 (p_0[28]), .A2 (Multiplier[28]));
NOR2_X1 slo__sro_c126 (.ZN (slo__sro_n195), .A1 (p_0[28]), .A2 (Multiplier[28]));
OAI21_X1 slo__sro_c127 (.ZN (slo__sro_n194), .A (slo__sro_n196), .B1 (slo__sro_n195), .B2 (slo__sro_n197));
NAND2_X1 slo__sro_c606 (.ZN (slo__sro_n882), .A1 (p_0[22]), .A2 (Multiplier[22]));
OAI21_X1 slo__sro_c607 (.ZN (slo__sro_n881), .A (slo__sro_n177), .B1 (p_0[22]), .B2 (Multiplier[22]));
NAND2_X1 slo__sro_c139 (.ZN (slo__sro_n212), .A1 (n_1), .A2 (Multiplier[1]));
NOR2_X1 slo__sro_c140 (.ZN (slo__sro_n211), .A1 (n_1), .A2 (Multiplier[1]));
OAI21_X1 slo__sro_c141 (.ZN (n_2), .A (slo__sro_n212), .B1 (slo__sro_n213), .B2 (slo__sro_n211));
XNOR2_X2 slo__sro_c142 (.ZN (slo__sro_n210), .A (n_1), .B (Multiplier[1]));
XNOR2_X1 slo__sro_c143 (.ZN (p_1[1]), .A (slo__sro_n210), .B (p_0[1]));
NAND2_X1 slo__sro_c153 (.ZN (slo__sro_n225), .A1 (n_7), .A2 (Multiplier[7]));
NOR2_X1 slo__sro_c154 (.ZN (slo__sro_n224), .A1 (n_7), .A2 (Multiplier[7]));
OAI21_X1 slo__sro_c155 (.ZN (n_8), .A (slo__sro_n225), .B1 (slo__sro_n226), .B2 (slo__sro_n224));
XNOR2_X2 slo__sro_c156 (.ZN (slo__sro_n223), .A (n_7), .B (Multiplier[7]));
XNOR2_X2 slo__sro_c157 (.ZN (p_1[7]), .A (slo__sro_n223), .B (p_0[7]));
NAND2_X1 slo__sro_c167 (.ZN (slo__sro_n241), .A1 (p_0[3]), .A2 (Multiplier[3]));
NOR2_X1 slo__sro_c168 (.ZN (slo__sro_n240), .A1 (p_0[3]), .A2 (Multiplier[3]));
OAI21_X1 slo__sro_c169 (.ZN (slo__sro_n239), .A (slo__sro_n241), .B1 (slo__sro_n242), .B2 (slo__sro_n240));
XNOR2_X2 slo__sro_c170 (.ZN (slo__sro_n238), .A (p_0[3]), .B (Multiplier[3]));
OR2_X1 CLOCK_slo__sro_c1214 (.ZN (CLOCK_slo__sro_n1759), .A1 (p_0[30]), .A2 (n_34));
NAND2_X1 slo__sro_c201 (.ZN (slo__sro_n280), .A1 (p_0[25]), .A2 (Multiplier[25]));
NOR2_X1 slo__sro_c202 (.ZN (slo__sro_n279), .A1 (p_0[25]), .A2 (Multiplier[25]));
OAI21_X1 slo__sro_c203 (.ZN (slo__sro_n278), .A (slo__sro_n280), .B1 (slo__sro_n279), .B2 (slo__sro_n281));
XNOR2_X2 slo__sro_c204 (.ZN (slo__sro_n277), .A (p_0[25]), .B (Multiplier[25]));
XNOR2_X2 slo__sro_c205 (.ZN (p_1[25]), .A (slo__sro_n277), .B (n_25));
INV_X1 slo__sro_c329 (.ZN (slo__sro_n464), .A (n_10));
NAND2_X1 slo__sro_c330 (.ZN (slo__sro_n463), .A1 (p_0[10]), .A2 (Multiplier[10]));
NOR2_X1 slo__sro_c331 (.ZN (slo__sro_n462), .A1 (p_0[10]), .A2 (Multiplier[10]));
OAI21_X1 slo__sro_c332 (.ZN (n_11), .A (slo__sro_n463), .B1 (slo__sro_n464), .B2 (slo__sro_n462));
XNOR2_X1 slo__sro_c333 (.ZN (slo__sro_n461), .A (p_0[10]), .B (Multiplier[10]));
INV_X1 slo__sro_c227 (.ZN (slo__sro_n309), .A (slo__sro_n647));
NAND2_X1 slo__sro_c228 (.ZN (slo__sro_n308), .A1 (p_0[17]), .A2 (Multiplier[17]));
NOR2_X1 slo__sro_c229 (.ZN (slo__sro_n307), .A1 (p_0[17]), .A2 (Multiplier[17]));
OAI21_X1 slo__sro_c230 (.ZN (n_18), .A (slo__sro_n308), .B1 (slo__sro_n309), .B2 (slo__sro_n307));
XNOR2_X2 slo__sro_c231 (.ZN (slo__sro_n306), .A (p_0[17]), .B (Multiplier[17]));
XNOR2_X1 slo__sro_c232 (.ZN (p_1[17]), .A (slo__sro_n306), .B (slo__sro_n647));
INV_X1 slo__sro_c401 (.ZN (slo__sro_n562), .A (n_27));
NOR2_X1 slo__sro_c403 (.ZN (slo__sro_n560), .A1 (p_0[27]), .A2 (Multiplier[27]));
OAI21_X4 slo__sro_c404 (.ZN (n_28), .A (slo__sro_n561), .B1 (slo__sro_n560), .B2 (slo__sro_n562));
XNOR2_X2 slo__sro_c405 (.ZN (slo__sro_n559), .A (p_0[27]), .B (Multiplier[27]));
XNOR2_X1 slo__sro_c406 (.ZN (p_1[27]), .A (slo__sro_n559), .B (n_27));
NAND2_X1 slo__sro_c464 (.ZN (slo__sro_n649), .A1 (p_0[16]), .A2 (Multiplier[16]));
NOR2_X1 slo__sro_c465 (.ZN (slo__sro_n648), .A1 (p_0[16]), .A2 (Multiplier[16]));
OAI21_X1 slo__sro_c466 (.ZN (slo__sro_n647), .A (slo__sro_n649), .B1 (slo__sro_n650), .B2 (slo__sro_n648));
XNOR2_X1 slo__sro_c467 (.ZN (slo__sro_n646), .A (p_0[16]), .B (Multiplier[16]));
XNOR2_X1 slo__sro_c468 (.ZN (p_1[16]), .A (slo__sro_n646), .B (n_16));
NAND2_X2 slo__sro_c608 (.ZN (n_23), .A1 (slo__sro_n881), .A2 (slo__sro_n882));
XNOR2_X1 slo__sro_c609 (.ZN (slo__sro_n880), .A (p_0[22]), .B (Multiplier[22]));
XNOR2_X1 slo__sro_c610 (.ZN (p_1[22]), .A (slo__sro_n880), .B (slo__sro_n177));
NAND2_X1 slo__sro_c627 (.ZN (slo__sro_n910), .A1 (opt_ipoPP_1), .A2 (Multiplier[9]));
NOR2_X1 slo__sro_c628 (.ZN (slo__sro_n909), .A1 (opt_ipoPP_1), .A2 (Multiplier[9]));
OAI21_X1 slo__sro_c629 (.ZN (n_10), .A (slo__sro_n910), .B1 (slo__sro_n911), .B2 (slo__sro_n909));
XNOR2_X1 slo__sro_c630 (.ZN (slo__sro_n908), .A (p_0[9]), .B (Multiplier[9]));
XNOR2_X1 slo__sro_c631 (.ZN (p_1[9]), .A (slo__sro_n908), .B (n_9));
NAND2_X1 CLOCK_slo__sro_c1010 (.ZN (CLOCK_slo__sro_n1525), .A1 (p_0[20]), .A2 (Multiplier[20]));
NOR2_X1 CLOCK_slo__sro_c1011 (.ZN (CLOCK_slo__sro_n1524), .A1 (p_0[20]), .A2 (Multiplier[20]));
NAND2_X1 CLOCK_slo__sro_c837 (.ZN (CLOCK_slo__sro_n1337), .A1 (p_0[5]), .A2 (Multiplier[5]));
OAI21_X2 CLOCK_slo__sro_c838 (.ZN (CLOCK_slo__sro_n1336), .A (n_5), .B1 (p_0[5]), .B2 (Multiplier[5]));
NAND2_X4 CLOCK_slo__sro_c839 (.ZN (n_6), .A1 (CLOCK_slo__sro_n1336), .A2 (CLOCK_slo__sro_n1337));
XNOR2_X2 CLOCK_slo__sro_c840 (.ZN (CLOCK_slo__sro_n1335), .A (p_0[5]), .B (Multiplier[5]));
XNOR2_X1 CLOCK_slo__sro_c841 (.ZN (p_1[5]), .A (CLOCK_slo__sro_n1335), .B (n_5));
XNOR2_X2 CLOCK_slo__mro_c897 (.ZN (p_1[6]), .A (CLOCK_slo__mro_n1383), .B (p_0[6]));
OAI21_X2 CLOCK_slo__sro_c1012 (.ZN (n_21), .A (CLOCK_slo__sro_n1525), .B1 (CLOCK_slo__sro_n1526), .B2 (CLOCK_slo__sro_n1524));
XNOR2_X1 CLOCK_slo__sro_c1013 (.ZN (CLOCK_slo__sro_n1523), .A (p_0[20]), .B (Multiplier[20]));
XNOR2_X1 CLOCK_slo__sro_c1014 (.ZN (p_1[20]), .A (CLOCK_slo__sro_n1523), .B (slo__sro_n88));

endmodule //datapath__0_196

module datapath__0_192 (opt_ipoPP_0, p_0, p_1, p_2);

output [31:0] p_2;
input [31:0] p_0;
input [31:0] p_1;
input opt_ipoPP_0;
wire spw_n1804;
wire slo__sro_n1097;
wire n_1;
wire n_2;
wire n_3;
wire n_4;
wire n_6;
wire n_7;
wire n_8;
wire n_9;
wire n_11;
wire n_12;
wire n_13;
wire n_15;
wire n_17;
wire n_19;
wire n_21;
wire n_22;
wire n_23;
wire n_24;
wire slo__sro_n1049;
wire n_26;
wire n_27;
wire n_28;
wire n_29;
wire n_30;
wire n_32;
wire n_0;
wire n_34;
wire n_33;
wire n_31;
wire slo__sro_n63;
wire slo__sro_n64;
wire slo__sro_n65;
wire slo__sro_n66;
wire slo__sro_n157;
wire slo__sro_n158;
wire slo__sro_n159;
wire slo__sro_n160;
wire slo__sro_n161;
wire CLOCK_slo__sro_n1543;
wire slo__sro_n175;
wire slo__sro_n176;
wire slo__sro_n177;
wire slo__sro_n178;
wire CLOCK_slo__sro_n1544;
wire CLOCK_slo__mro_n1533;
wire slo__sro_n388;
wire slo__sro_n389;
wire CLOCK_slo__sro_n1561;
wire slo__sro_n221;
wire slo__sro_n222;
wire slo__sro_n223;
wire slo__sro_n224;
wire CLOCK_slo__sro_n1560;
wire slo__sro_n350;
wire slo__sro_n351;
wire slo__sro_n352;
wire slo__sro_n390;
wire slo__sro_n443;
wire slo__sro_n444;
wire slo__sro_n445;
wire slo__sro_n446;
wire slo__sro_n447;
wire slo__sro_n535;
wire slo__sro_n536;
wire slo__sro_n537;
wire slo__sro_n538;
wire slo__sro_n550;
wire slo__sro_n551;
wire slo__sro_n552;
wire slo__sro_n553;
wire slo__sro_n703;
wire slo__sro_n704;
wire slo__sro_n705;
wire slo__sro_n706;
wire slo__sro_n995;
wire slo__sro_n996;
wire slo__sro_n997;
wire slo__sro_n998;
wire slo__sro_n1093;
wire slo__sro_n1094;
wire slo__sro_n1095;
wire slo__sro_n1096;
wire slo__sro_n1045;
wire slo__sro_n1046;
wire slo__sro_n1047;
wire slo__sro_n1048;
wire slo__sro_n759;
wire slo__sro_n760;
wire slo__sro_n761;
wire slo__sro_n762;
wire slo__sro_n763;
wire slo__sro_n1050;
wire CLOCK_slo__mro_n1516;
wire CLOCK_slo__sro_n1545;
wire CLOCK_slo__mro_n1551;
wire CLOCK_slo__sro_n1562;
wire CLOCK_slo__sro_n1563;
wire CLOCK_slo__sro_n1570;
wire CLOCK_slo__sro_n1571;
wire CLOCK_slo__sro_n1572;
wire CLOCK_slo__sro_n1573;
wire slo__sro_n1427;
wire slo__sro_n1429;
wire CLOCK_slo__sro_n1719;
wire CLOCK_slo__sro_n1720;
wire CLOCK_slo__sro_n1721;
wire CLOCK_slo__sro_n1722;


INV_X1 i_36 (.ZN (n_34), .A (p_0[30]));
INV_X1 i_35 (.ZN (n_33), .A (p_1[30]));
INV_X1 i_34 (.ZN (n_32), .A (n_30));
INV_X1 CLOCK_slo__sro_c1046 (.ZN (CLOCK_slo__sro_n1573), .A (p_1[20]));
XOR2_X1 i_32 (.Z (p_2[31]), .A (p_0[31]), .B (n_31));
OAI22_X1 i_31 (.ZN (n_0), .A1 (n_34), .A2 (p_1[30]), .B1 (p_0[30]), .B2 (n_33));
XNOR2_X1 i_0 (.ZN (p_2[30]), .A (n_32), .B (n_0));
FA_X1 i_30 (.CO (n_30), .S (p_2[29]), .A (p_0[29]), .B (spw_n1804), .CI (n_29));
FA_X1 i_29 (.CO (n_29), .S (p_2[28]), .A (p_0[28]), .B (p_1[28]), .CI (n_28));
INV_X1 slo__sro_c774 (.ZN (slo__sro_n1097), .A (n_17));
FA_X1 i_27 (.CO (n_27), .S (p_2[26]), .A (p_0[26]), .B (p_1[26]), .CI (n_26));
XNOR2_X2 CLOCK_slo__mro_c987 (.ZN (p_2[3]), .A (CLOCK_slo__mro_n1516), .B (n_3));
XNOR2_X1 slo__sro_c752 (.ZN (slo__sro_n1045), .A (p_1[25]), .B (p_0[25]));
FA_X1 i_24 (.CO (n_24), .S (p_2[23]), .A (p_0[23]), .B (p_1[23]), .CI (n_23));
FA_X1 i_23 (.CO (n_23), .S (p_2[22]), .A (p_0[22]), .B (p_1[22]), .CI (n_22));
FA_X1 i_22 (.CO (n_22), .S (p_2[21]), .A (p_0[21]), .B (p_1[21]), .CI (n_21));
INV_X1 CLOCK_slo__sro_c1151 (.ZN (CLOCK_slo__sro_n1722), .A (n_6));
XNOR2_X1 CLOCK_slo__mro_c1024 (.ZN (CLOCK_slo__mro_n1551), .A (p_1[7]), .B (p_0[7]));
FA_X1 i_19 (.CO (n_19), .S (p_2[18]), .A (p_0[18]), .B (p_1[18]), .CI (slo__sro_n1094));
XNOR2_X2 CLOCK_slo__mro_c986 (.ZN (CLOCK_slo__mro_n1516), .A (p_1[3]), .B (p_0[3]));
FA_X1 i_17 (.CO (n_17), .S (p_2[16]), .A (p_0[16]), .B (p_1[16]), .CI (slo__sro_n704));
NAND2_X1 slo__sro_c709 (.ZN (slo__sro_n997), .A1 (p_1[27]), .A2 (p_0[27]));
INV_X1 slo__sro_c271 (.ZN (slo__sro_n352), .A (n_7));
INV_X1 slo__sro_c107 (.ZN (slo__sro_n178), .A (n_19));
FA_X1 i_13 (.CO (n_13), .S (p_2[12]), .A (p_0[12]), .B (p_1[12]), .CI (n_12));
FA_X1 i_12 (.CO (n_12), .S (p_2[11]), .A (p_0[11]), .B (p_1[11]), .CI (n_11));
INV_X1 slo__sro_c93 (.ZN (slo__sro_n161), .A (n_13));
NAND2_X1 slo__sro_c402 (.ZN (slo__sro_n553), .A1 (opt_ipoPP_0), .A2 (p_0[4]));
FA_X1 i_9 (.CO (n_9), .S (p_2[8]), .A (p_0[8]), .B (p_1[8]), .CI (n_8));
INV_X1 CLOCK_slo__sro_c1015 (.ZN (CLOCK_slo__sro_n1544), .A (p_0[15]));
FA_X1 i_6 (.CO (n_6), .S (p_2[5]), .A (p_0[5]), .B (p_1[5]), .CI (slo__sro_n551));
INV_X1 slo__sro_c708 (.ZN (slo__sro_n998), .A (n_27));
INV_X1 slo__sro_c324 (.ZN (slo__sro_n447), .A (n_9));
XNOR2_X1 CLOCK_slo__mro_c1004 (.ZN (CLOCK_slo__mro_n1533), .A (p_1[19]), .B (p_0[19]));
FA_X1 i_2 (.CO (n_2), .S (p_2[1]), .A (p_0[1]), .B (p_1[1]), .CI (n_1));
HA_X1 i_1 (.CO (n_1), .S (p_2[0]), .A (p_0[0]), .B (p_1[0]));
INV_X1 slo__sro_c1 (.ZN (slo__sro_n66), .A (slo__sro_n444));
NAND2_X1 slo__sro_c2 (.ZN (slo__sro_n65), .A1 (p_1[10]), .A2 (p_0[10]));
NOR2_X1 slo__sro_c3 (.ZN (slo__sro_n64), .A1 (p_1[10]), .A2 (p_0[10]));
OAI21_X1 slo__sro_c4 (.ZN (n_11), .A (slo__sro_n65), .B1 (slo__sro_n66), .B2 (slo__sro_n64));
XNOR2_X1 slo__sro_c5 (.ZN (slo__sro_n63), .A (p_1[10]), .B (p_0[10]));
XNOR2_X1 slo__sro_c6 (.ZN (p_2[10]), .A (slo__sro_n63), .B (slo__sro_n444));
NAND2_X1 slo__sro_c94 (.ZN (slo__sro_n160), .A1 (p_1[13]), .A2 (p_0[13]));
NOR2_X1 slo__sro_c95 (.ZN (slo__sro_n159), .A1 (p_1[13]), .A2 (p_0[13]));
OAI21_X2 slo__sro_c96 (.ZN (slo__sro_n158), .A (slo__sro_n160), .B1 (slo__sro_n161), .B2 (slo__sro_n159));
XNOR2_X1 slo__sro_c97 (.ZN (slo__sro_n157), .A (p_1[13]), .B (p_0[13]));
XNOR2_X1 slo__sro_c98 (.ZN (p_2[13]), .A (slo__sro_n157), .B (n_13));
NAND2_X1 slo__sro_c108 (.ZN (slo__sro_n177), .A1 (p_1[19]), .A2 (p_0[19]));
NOR2_X1 slo__sro_c109 (.ZN (slo__sro_n176), .A1 (p_1[19]), .A2 (p_0[19]));
OAI21_X1 slo__sro_c110 (.ZN (slo__sro_n175), .A (slo__sro_n177), .B1 (slo__sro_n178), .B2 (slo__sro_n176));
INV_X1 CLOCK_slo__sro_c1014 (.ZN (CLOCK_slo__sro_n1545), .A (p_1[15]));
XNOR2_X1 slo__sro_c112 (.ZN (p_2[19]), .A (CLOCK_slo__mro_n1533), .B (n_19));
INV_X2 slo__sro_c296 (.ZN (slo__sro_n390), .A (n_3));
NAND2_X1 slo__sro_c297 (.ZN (slo__sro_n389), .A1 (p_0[3]), .A2 (p_1[3]));
NOR2_X1 slo__sro_c298 (.ZN (slo__sro_n388), .A1 (p_1[3]), .A2 (p_0[3]));
OAI21_X1 slo__sro_c299 (.ZN (n_4), .A (slo__sro_n389), .B1 (slo__sro_n388), .B2 (slo__sro_n390));
OAI21_X1 CLOCK_slo__sro_c1000 (.ZN (slo__sro_n552), .A (n_4), .B1 (p_1[4]), .B2 (p_0[4]));
INV_X1 slo__sro_c147 (.ZN (slo__sro_n224), .A (p_1[14]));
NAND2_X1 slo__sro_c148 (.ZN (slo__sro_n223), .A1 (slo__sro_n158), .A2 (p_0[14]));
NOR2_X1 slo__sro_c149 (.ZN (slo__sro_n222), .A1 (slo__sro_n158), .A2 (p_0[14]));
OAI21_X1 slo__sro_c150 (.ZN (n_15), .A (slo__sro_n223), .B1 (slo__sro_n224), .B2 (slo__sro_n222));
XNOR2_X1 slo__sro_c151 (.ZN (slo__sro_n221), .A (slo__sro_n158), .B (p_0[14]));
XNOR2_X1 slo__sro_c152 (.ZN (p_2[14]), .A (slo__sro_n221), .B (p_1[14]));
NAND2_X1 slo__sro_c272 (.ZN (slo__sro_n351), .A1 (p_1[7]), .A2 (p_0[7]));
NOR2_X1 slo__sro_c273 (.ZN (slo__sro_n350), .A1 (p_1[7]), .A2 (p_0[7]));
OAI21_X1 slo__sro_c274 (.ZN (n_8), .A (slo__sro_n351), .B1 (slo__sro_n352), .B2 (slo__sro_n350));
INV_X1 CLOCK_slo__sro_c1032 (.ZN (CLOCK_slo__sro_n1563), .A (n_30));
NOR2_X1 CLOCK_slo__sro_c1033 (.ZN (CLOCK_slo__sro_n1562), .A1 (n_33), .A2 (p_0[30]));
NAND2_X1 slo__sro_c325 (.ZN (slo__sro_n446), .A1 (p_1[9]), .A2 (p_0[9]));
NOR2_X1 slo__sro_c326 (.ZN (slo__sro_n445), .A1 (p_1[9]), .A2 (p_0[9]));
OAI21_X1 slo__sro_c327 (.ZN (slo__sro_n444), .A (slo__sro_n446), .B1 (slo__sro_n447), .B2 (slo__sro_n445));
XNOR2_X2 slo__sro_c328 (.ZN (slo__sro_n443), .A (p_1[9]), .B (p_0[9]));
XNOR2_X1 slo__sro_c329 (.ZN (p_2[9]), .A (slo__sro_n443), .B (n_9));
INV_X1 slo__sro_c386 (.ZN (slo__sro_n538), .A (n_2));
NAND2_X1 slo__sro_c387 (.ZN (slo__sro_n537), .A1 (p_1[2]), .A2 (p_0[2]));
NOR2_X1 slo__sro_c388 (.ZN (slo__sro_n536), .A1 (p_1[2]), .A2 (p_0[2]));
OAI21_X2 slo__sro_c389 (.ZN (n_3), .A (slo__sro_n537), .B1 (slo__sro_n536), .B2 (slo__sro_n538));
XNOR2_X1 slo__sro_c390 (.ZN (slo__sro_n535), .A (p_1[2]), .B (p_0[2]));
XNOR2_X1 slo__sro_c391 (.ZN (p_2[2]), .A (slo__sro_n535), .B (n_2));
NAND2_X1 slo__sro_c404 (.ZN (slo__sro_n551), .A1 (slo__sro_n552), .A2 (slo__sro_n553));
XNOR2_X1 slo__sro_c405 (.ZN (slo__sro_n550), .A (n_4), .B (p_0[4]));
XNOR2_X1 slo__sro_c406 (.ZN (p_2[4]), .A (slo__sro_n550), .B (opt_ipoPP_0));
NAND2_X1 slo__sro_c508 (.ZN (slo__sro_n706), .A1 (p_1[15]), .A2 (p_0[15]));
NAND2_X1 slo__sro_c510 (.ZN (slo__sro_n704), .A1 (slo__sro_n705), .A2 (slo__sro_n706));
XNOR2_X1 slo__sro_c511 (.ZN (slo__sro_n703), .A (p_1[15]), .B (p_0[15]));
XNOR2_X1 slo__sro_c512 (.ZN (p_2[15]), .A (slo__sro_n703), .B (n_15));
NOR2_X1 slo__sro_c710 (.ZN (slo__sro_n996), .A1 (p_1[27]), .A2 (p_0[27]));
OAI21_X1 slo__sro_c711 (.ZN (n_28), .A (slo__sro_n997), .B1 (slo__sro_n998), .B2 (slo__sro_n996));
XNOR2_X1 slo__sro_c712 (.ZN (slo__sro_n995), .A (p_1[27]), .B (p_0[27]));
XNOR2_X1 slo__sro_c713 (.ZN (p_2[27]), .A (slo__sro_n995), .B (n_27));
NAND2_X1 slo__sro_c775 (.ZN (slo__sro_n1096), .A1 (p_1[17]), .A2 (p_0[17]));
NOR2_X1 slo__sro_c776 (.ZN (slo__sro_n1095), .A1 (p_1[17]), .A2 (p_0[17]));
OAI21_X1 slo__sro_c777 (.ZN (slo__sro_n1094), .A (slo__sro_n1096), .B1 (slo__sro_n1097), .B2 (slo__sro_n1095));
XNOR2_X1 slo__sro_c778 (.ZN (slo__sro_n1093), .A (p_1[17]), .B (p_0[17]));
XNOR2_X1 slo__sro_c779 (.ZN (p_2[17]), .A (slo__sro_n1093), .B (n_17));
INV_X1 slo__sro_c746 (.ZN (slo__sro_n1050), .A (p_0[25]));
INV_X1 slo__sro_c747 (.ZN (slo__sro_n1049), .A (p_1[25]));
NAND2_X1 slo__sro_c748 (.ZN (slo__sro_n1048), .A1 (p_1[25]), .A2 (p_0[25]));
NAND2_X1 slo__sro_c749 (.ZN (slo__sro_n1047), .A1 (slo__sro_n1050), .A2 (slo__sro_n1049));
NAND2_X1 slo__sro_c750 (.ZN (slo__sro_n1046), .A1 (slo__sro_n760), .A2 (slo__sro_n1047));
NAND2_X1 slo__sro_c751 (.ZN (n_26), .A1 (slo__sro_n1048), .A2 (slo__sro_n1046));
INV_X1 slo__sro_c559 (.ZN (slo__sro_n763), .A (n_24));
NAND2_X1 slo__sro_c560 (.ZN (slo__sro_n762), .A1 (p_1[24]), .A2 (p_0[24]));
NOR2_X1 slo__sro_c561 (.ZN (slo__sro_n761), .A1 (p_1[24]), .A2 (p_0[24]));
OAI21_X2 slo__sro_c562 (.ZN (slo__sro_n760), .A (slo__sro_n762), .B1 (slo__sro_n763), .B2 (slo__sro_n761));
XNOR2_X1 slo__sro_c563 (.ZN (slo__sro_n759), .A (p_1[24]), .B (p_0[24]));
XNOR2_X1 slo__sro_c564 (.ZN (p_2[24]), .A (n_24), .B (slo__sro_n759));
XNOR2_X2 slo__sro_c753 (.ZN (p_2[25]), .A (slo__sro_n1045), .B (slo__sro_n760));
NAND2_X1 CLOCK_slo__sro_c1016 (.ZN (CLOCK_slo__sro_n1543), .A1 (CLOCK_slo__sro_n1544), .A2 (CLOCK_slo__sro_n1545));
NAND2_X1 CLOCK_slo__sro_c1017 (.ZN (slo__sro_n705), .A1 (CLOCK_slo__sro_n1543), .A2 (n_15));
XNOR2_X1 CLOCK_slo__mro_c1025 (.ZN (p_2[7]), .A (CLOCK_slo__mro_n1551), .B (n_7));
NAND2_X1 CLOCK_slo__sro_c1034 (.ZN (CLOCK_slo__sro_n1561), .A1 (CLOCK_slo__sro_n1563), .A2 (CLOCK_slo__sro_n1562));
OR2_X1 CLOCK_slo__sro_c1035 (.ZN (CLOCK_slo__sro_n1560), .A1 (p_1[30]), .A2 (n_34));
OAI21_X1 CLOCK_slo__sro_c1036 (.ZN (n_31), .A (CLOCK_slo__sro_n1561), .B1 (n_32), .B2 (CLOCK_slo__sro_n1560));
INV_X1 CLOCK_slo__sro_c1047 (.ZN (CLOCK_slo__sro_n1572), .A (p_0[20]));
NAND2_X1 CLOCK_slo__sro_c1048 (.ZN (CLOCK_slo__sro_n1571), .A1 (CLOCK_slo__sro_n1572), .A2 (CLOCK_slo__sro_n1573));
NAND2_X1 CLOCK_slo__sro_c1049 (.ZN (CLOCK_slo__sro_n1570), .A1 (CLOCK_slo__sro_n1571), .A2 (slo__sro_n175));
CLKBUF_X1 spw__L1_c1_c1242 (.Z (spw_n1804), .A (p_1[29]));
NAND2_X1 slo__sro_c941 (.ZN (slo__sro_n1429), .A1 (p_1[20]), .A2 (p_0[20]));
NAND2_X1 slo__sro_c943 (.ZN (n_21), .A1 (slo__sro_n1429), .A2 (CLOCK_slo__sro_n1570));
XNOR2_X1 slo__sro_c944 (.ZN (slo__sro_n1427), .A (p_1[20]), .B (p_0[20]));
XNOR2_X1 slo__sro_c945 (.ZN (p_2[20]), .A (slo__sro_n1427), .B (slo__sro_n175));
NAND2_X1 CLOCK_slo__sro_c1152 (.ZN (CLOCK_slo__sro_n1721), .A1 (p_1[6]), .A2 (p_0[6]));
NOR2_X1 CLOCK_slo__sro_c1153 (.ZN (CLOCK_slo__sro_n1720), .A1 (p_1[6]), .A2 (p_0[6]));
OAI21_X2 CLOCK_slo__sro_c1154 (.ZN (n_7), .A (CLOCK_slo__sro_n1721), .B1 (CLOCK_slo__sro_n1722), .B2 (CLOCK_slo__sro_n1720));
XNOR2_X1 CLOCK_slo__sro_c1155 (.ZN (CLOCK_slo__sro_n1719), .A (p_1[6]), .B (p_0[6]));
XNOR2_X1 CLOCK_slo__sro_c1156 (.ZN (p_2[6]), .A (CLOCK_slo__sro_n1719), .B (n_6));

endmodule //datapath__0_192

module datapath__0_191 (Multiplier, p_0, p_1);

output [31:0] p_1;
input [31:0] Multiplier;
input [31:0] p_0;
wire CLOCK_slo__sro_n1159;
wire slo__sro_n550;
wire n_1;
wire n_2;
wire n_3;
wire n_4;
wire n_5;
wire n_6;
wire n_7;
wire n_8;
wire n_10;
wire n_11;
wire n_12;
wire n_13;
wire n_14;
wire n_15;
wire n_16;
wire n_17;
wire slo__sro_n877;
wire n_19;
wire n_23;
wire n_25;
wire n_26;
wire n_28;
wire n_30;
wire n_32;
wire CLOCK_slo__sro_n1408;
wire n_34;
wire n_33;
wire slo__sro_n57;
wire slo__sro_n58;
wire slo__sro_n59;
wire slo__sro_n60;
wire slo__sro_n813;
wire slo__sro_n71;
wire slo__sro_n72;
wire slo__sro_n73;
wire slo__sro_n74;
wire slo__sro_n87;
wire slo__sro_n88;
wire slo__sro_n89;
wire slo__sro_n90;
wire slo__sro_n100;
wire slo__sro_n101;
wire slo__sro_n102;
wire slo__sro_n103;
wire slo__sro_n128;
wire slo__sro_n129;
wire slo__sro_n130;
wire slo__sro_n131;
wire slo__sro_n141;
wire slo__sro_n142;
wire slo__sro_n143;
wire slo__sro_n144;
wire slo__sro_n156;
wire slo__sro_n157;
wire slo__sro_n158;
wire slo__sro_n159;
wire slo__sro_n175;
wire slo__sro_n176;
wire slo__sro_n185;
wire slo__sro_n186;
wire slo__sro_n187;
wire slo__sro_n188;
wire slo__sro_n189;
wire CLOCK_slo__sro_n1158;
wire slo__sro_n205;
wire slo__sro_n206;
wire slo__sro_n293;
wire slo__n250;
wire CLOCK_slo__sro_n1192;
wire slo__sro_n295;
wire slo__sro_n296;
wire slo__sro_n325;
wire slo__sro_n326;
wire slo__sro_n327;
wire slo__sro_n328;
wire slo__sro_n329;
wire slo__sro_n551;
wire slo__sro_n552;
wire slo__sro_n553;
wire slo__sro_n741;
wire slo__sro_n742;
wire slo__xsl_n702;
wire slo__xsl_n703;
wire slo__sro_n739;
wire slo__sro_n740;
wire slo__mro_n781;
wire slo__sro_n814;
wire slo__sro_n815;
wire slo__sro_n816;
wire slo__mro_n862;
wire slo__sro_n878;
wire slo__sro_n879;
wire slo__sro_n880;
wire CLOCK_slo__mro_n1145;
wire CLOCK_slo__sro_n1160;
wire CLOCK_slo__sro_n1161;
wire CLOCK_slo__sro_n1162;
wire CLOCK_slo__mro_n1184;
wire CLOCK_slo__sro_n1193;
wire CLOCK_slo__sro_n1194;
wire CLOCK_slo__sro_n1195;
wire CLOCK_slo__sro_n1223;
wire CLOCK_slo__sro_n1224;
wire CLOCK_slo__sro_n1225;
wire CLOCK_slo__sro_n1226;
wire CLOCK_slo__sro_n1250;
wire CLOCK_slo__sro_n1251;
wire CLOCK_slo__sro_n1252;
wire CLOCK_slo__sro_n1253;
wire CLOCK_slo__sro_n1254;
wire CLOCK_slo__sro_n1269;
wire CLOCK_slo__sro_n1270;
wire CLOCK_slo__sro_n1271;
wire CLOCK_slo__sro_n1272;
wire CLOCK_slo__sro_n1294;
wire CLOCK_slo__sro_n1409;
wire CLOCK_slo__sro_n1410;
wire CLOCK_slo__sro_n1411;


INV_X1 i_36 (.ZN (n_34), .A (Multiplier[30]));
INV_X2 i_35 (.ZN (n_33), .A (p_0[30]));
INV_X1 i_34 (.ZN (n_32), .A (n_30));
INV_X1 CLOCK_slo__sro_c787 (.ZN (CLOCK_slo__sro_n1195), .A (CLOCK_slo__sro_n1270));
XOR2_X1 i_32 (.Z (p_1[31]), .A (Multiplier[31]), .B (CLOCK_slo__sro_n1158));
NAND2_X1 CLOCK_slo__sro_c928 (.ZN (CLOCK_slo__sro_n1410), .A1 (n_2), .A2 (Multiplier[2]));
XNOR2_X1 i_0 (.ZN (p_1[30]), .A (n_32), .B (CLOCK_slo__sro_n1294));
FA_X1 i_30 (.CO (n_30), .S (p_1[29]), .A (Multiplier[29]), .B (p_0[29]), .CI (CLOCK_slo__sro_n1224));
INV_X1 CLOCK_slo__sro_c838 (.ZN (CLOCK_slo__sro_n1254), .A (n_8));
XNOR2_X1 slo__mro_c596 (.ZN (slo__mro_n862), .A (p_0[15]), .B (Multiplier[15]));
NAND2_X1 slo__sro_c141 (.ZN (slo__sro_n206), .A1 (p_0[4]), .A2 (Multiplier[4]));
FA_X1 i_26 (.CO (n_26), .S (p_1[25]), .A (Multiplier[25]), .B (p_0[25]), .CI (n_25));
NAND2_X1 slo__sro_c86 (.ZN (slo__sro_n144), .A1 (slo__sro_n71), .A2 (Multiplier[20]));
NAND2_X1 slo__sro_c372 (.ZN (slo__sro_n552), .A1 (p_0[9]), .A2 (Multiplier[9]));
NAND2_X1 CLOCK_slo__sro_c813 (.ZN (CLOCK_slo__sro_n1226), .A1 (p_0[28]), .A2 (Multiplier[28]));
NAND2_X1 CLOCK_slo__sro_c927 (.ZN (CLOCK_slo__sro_n1411), .A1 (p_0[2]), .A2 (Multiplier[2]));
NAND2_X1 slo__sro_c98 (.ZN (slo__sro_n159), .A1 (p_0[17]), .A2 (Multiplier[17]));
INV_X1 slo__sro_c29 (.ZN (slo__sro_n90), .A (n_5));
XNOR2_X2 CLOCK_slo__mro_c735 (.ZN (CLOCK_slo__mro_n1145), .A (p_0[4]), .B (Multiplier[4]));
NAND2_X1 slo__sro_c113 (.ZN (slo__sro_n176), .A1 (n_15), .A2 (Multiplier[15]));
FA_X1 i_17 (.CO (n_17), .S (p_1[16]), .A (Multiplier[16]), .B (p_0[16]), .CI (n_16));
INV_X1 slo__sro_c125 (.ZN (slo__sro_n189), .A (n_26));
INV_X1 slo__sro_c72 (.ZN (slo__sro_n131), .A (slo__sro_n326));
FA_X1 i_14 (.CO (n_14), .S (p_1[13]), .A (Multiplier[13]), .B (p_0[13]), .CI (n_13));
INV_X1 slo__sro_c15 (.ZN (slo__sro_n74), .A (n_19));
XNOR2_X2 slo__mro_c531 (.ZN (slo__mro_n781), .A (p_0[19]), .B (Multiplier[19]));
FA_X1 i_11 (.CO (n_11), .S (p_1[10]), .A (Multiplier[10]), .B (p_0[10]), .CI (n_10));
XNOR2_X1 slo__sro_c506 (.ZN (slo__sro_n739), .A (p_0[11]), .B (Multiplier[11]));
NAND2_X1 CLOCK_slo__sro_c854 (.ZN (CLOCK_slo__sro_n1272), .A1 (p_0[21]), .A2 (Multiplier[21]));
FA_X1 i_8 (.CO (n_8), .S (p_1[7]), .A (Multiplier[7]), .B (p_0[7]), .CI (n_7));
FA_X1 i_7 (.CO (n_7), .S (p_1[6]), .A (Multiplier[6]), .B (p_0[6]), .CI (n_6));
INV_X1 slo__sro_c43 (.ZN (slo__sro_n103), .A (n_14));
INV_X1 slo__sro_c371 (.ZN (slo__sro_n553), .A (CLOCK_slo__sro_n1251));
INV_X1 slo__sro_c226 (.ZN (slo__sro_n329), .A (n_23));
FA_X1 i_2 (.CO (n_2), .S (p_1[1]), .A (Multiplier[1]), .B (p_0[1]), .CI (n_1));
HA_X1 i_1 (.CO (n_1), .S (p_1[0]), .A (Multiplier[0]), .B (p_0[0]));
INV_X1 slo__sro_c1 (.ZN (slo__sro_n60), .A (n_12));
NAND2_X1 slo__sro_c2 (.ZN (slo__sro_n59), .A1 (p_0[12]), .A2 (Multiplier[12]));
NOR2_X1 slo__sro_c3 (.ZN (slo__sro_n58), .A1 (p_0[12]), .A2 (Multiplier[12]));
OAI21_X1 slo__sro_c4 (.ZN (n_13), .A (slo__sro_n59), .B1 (slo__sro_n60), .B2 (slo__sro_n58));
XNOR2_X1 slo__sro_c5 (.ZN (slo__sro_n57), .A (p_0[12]), .B (Multiplier[12]));
INV_X1 slo__sro_c502 (.ZN (slo__sro_n742), .A (n_11));
NAND2_X1 slo__sro_c16 (.ZN (slo__sro_n73), .A1 (p_0[19]), .A2 (Multiplier[19]));
NOR2_X1 slo__sro_c17 (.ZN (slo__sro_n72), .A1 (p_0[19]), .A2 (Multiplier[19]));
OAI21_X1 slo__sro_c18 (.ZN (slo__sro_n71), .A (slo__sro_n73), .B1 (slo__sro_n72), .B2 (slo__sro_n74));
INV_X1 slo__sro_c549 (.ZN (slo__sro_n816), .A (p_0[27]));
NAND2_X1 slo__sro_c550 (.ZN (slo__sro_n815), .A1 (slo__sro_n186), .A2 (Multiplier[27]));
NAND2_X1 slo__sro_c30 (.ZN (slo__sro_n89), .A1 (p_0[5]), .A2 (Multiplier[5]));
NOR2_X1 slo__sro_c31 (.ZN (slo__sro_n88), .A1 (p_0[5]), .A2 (Multiplier[5]));
OAI21_X2 slo__sro_c32 (.ZN (n_6), .A (slo__sro_n89), .B1 (slo__sro_n88), .B2 (slo__sro_n90));
XNOR2_X1 slo__sro_c33 (.ZN (slo__sro_n87), .A (p_0[5]), .B (Multiplier[5]));
XNOR2_X1 slo__sro_c34 (.ZN (p_1[5]), .A (slo__sro_n87), .B (n_5));
NAND2_X1 slo__sro_c44 (.ZN (slo__sro_n102), .A1 (p_0[14]), .A2 (Multiplier[14]));
NOR2_X1 slo__sro_c608 (.ZN (slo__sro_n878), .A1 (p_0[18]), .A2 (Multiplier[18]));
OAI21_X1 slo__sro_c46 (.ZN (n_15), .A (slo__sro_n102), .B1 (slo__sro_n103), .B2 (slo__sro_n101));
XNOR2_X1 slo__sro_c47 (.ZN (slo__sro_n100), .A (p_0[14]), .B (Multiplier[14]));
XNOR2_X1 slo__sro_c48 (.ZN (p_1[14]), .A (slo__sro_n100), .B (n_14));
NAND2_X1 slo__sro_c73 (.ZN (slo__sro_n130), .A1 (p_0[24]), .A2 (Multiplier[24]));
NOR2_X1 slo__sro_c74 (.ZN (slo__sro_n129), .A1 (p_0[24]), .A2 (Multiplier[24]));
OAI21_X1 slo__sro_c75 (.ZN (n_25), .A (slo__sro_n130), .B1 (slo__sro_n129), .B2 (slo__sro_n131));
XNOR2_X2 slo__sro_c76 (.ZN (slo__sro_n128), .A (p_0[24]), .B (Multiplier[24]));
XNOR2_X2 slo__sro_c77 (.ZN (p_1[24]), .A (slo__sro_n128), .B (slo__xsl_n702));
OAI21_X1 slo__sro_c87 (.ZN (slo__sro_n143), .A (p_0[20]), .B1 (slo__sro_n71), .B2 (Multiplier[20]));
NAND2_X1 slo__sro_c88 (.ZN (slo__sro_n142), .A1 (slo__sro_n143), .A2 (slo__sro_n144));
XNOR2_X1 slo__sro_c89 (.ZN (slo__sro_n141), .A (slo__sro_n71), .B (Multiplier[20]));
XNOR2_X1 slo__sro_c90 (.ZN (p_1[20]), .A (slo__sro_n141), .B (p_0[20]));
OAI21_X1 slo__sro_c99 (.ZN (slo__sro_n158), .A (n_17), .B1 (p_0[17]), .B2 (Multiplier[17]));
NAND2_X1 slo__sro_c100 (.ZN (slo__sro_n157), .A1 (slo__sro_n159), .A2 (slo__sro_n158));
XNOR2_X1 slo__sro_c101 (.ZN (slo__sro_n156), .A (p_0[17]), .B (Multiplier[17]));
XNOR2_X1 slo__sro_c102 (.ZN (p_1[17]), .A (slo__sro_n156), .B (n_17));
OAI21_X1 slo__sro_c114 (.ZN (slo__sro_n175), .A (p_0[15]), .B1 (slo__n250), .B2 (Multiplier[15]));
NAND2_X1 slo__sro_c115 (.ZN (n_16), .A1 (slo__sro_n175), .A2 (slo__sro_n176));
INV_X1 slo__sro_c606 (.ZN (slo__sro_n880), .A (slo__sro_n157));
NAND2_X1 slo__sro_c607 (.ZN (slo__sro_n879), .A1 (p_0[18]), .A2 (Multiplier[18]));
NAND2_X1 slo__sro_c126 (.ZN (slo__sro_n188), .A1 (p_0[26]), .A2 (Multiplier[26]));
NOR2_X1 slo__sro_c127 (.ZN (slo__sro_n187), .A1 (p_0[26]), .A2 (Multiplier[26]));
OAI21_X2 slo__sro_c128 (.ZN (slo__sro_n186), .A (slo__sro_n188), .B1 (slo__sro_n187), .B2 (slo__sro_n189));
XNOR2_X2 slo__sro_c129 (.ZN (slo__sro_n185), .A (p_0[26]), .B (Multiplier[26]));
XNOR2_X2 slo__sro_c130 (.ZN (p_1[26]), .A (slo__sro_n185), .B (n_26));
OAI21_X1 slo__sro_c142 (.ZN (slo__sro_n205), .A (n_4), .B1 (p_0[4]), .B2 (Multiplier[4]));
NAND2_X2 slo__sro_c143 (.ZN (n_5), .A1 (slo__sro_n206), .A2 (slo__sro_n205));
INV_X1 CLOCK_slo__sro_c747 (.ZN (CLOCK_slo__sro_n1162), .A (n_30));
NOR2_X1 CLOCK_slo__sro_c748 (.ZN (CLOCK_slo__sro_n1161), .A1 (n_33), .A2 (Multiplier[30]));
INV_X1 slo__sro_c202 (.ZN (slo__sro_n296), .A (n_3));
NAND2_X1 slo__sro_c203 (.ZN (slo__sro_n295), .A1 (p_0[3]), .A2 (Multiplier[3]));
OAI21_X1 slo__c178 (.ZN (slo__n250), .A (slo__sro_n102), .B1 (slo__sro_n103), .B2 (slo__sro_n101));
NOR2_X1 CLOCK_slo__sro_c789 (.ZN (CLOCK_slo__sro_n1193), .A1 (p_0[22]), .A2 (Multiplier[22]));
OAI21_X2 slo__sro_c205 (.ZN (n_4), .A (slo__sro_n295), .B1 (CLOCK_slo__mro_n1184), .B2 (slo__sro_n296));
XNOR2_X1 slo__sro_c206 (.ZN (slo__sro_n293), .A (p_0[3]), .B (Multiplier[3]));
XNOR2_X1 slo__sro_c207 (.ZN (p_1[3]), .A (slo__sro_n293), .B (n_3));
NAND2_X1 slo__sro_c227 (.ZN (slo__sro_n328), .A1 (p_0[23]), .A2 (Multiplier[23]));
NOR2_X1 slo__sro_c228 (.ZN (slo__sro_n327), .A1 (p_0[23]), .A2 (Multiplier[23]));
OAI21_X2 slo__sro_c229 (.ZN (slo__sro_n326), .A (slo__sro_n328), .B1 (slo__sro_n329), .B2 (slo__sro_n327));
XNOR2_X1 slo__sro_c230 (.ZN (slo__sro_n325), .A (p_0[23]), .B (Multiplier[23]));
XNOR2_X1 slo__sro_c231 (.ZN (p_1[23]), .A (slo__sro_n325), .B (n_23));
NOR2_X1 slo__sro_c373 (.ZN (slo__sro_n551), .A1 (p_0[9]), .A2 (Multiplier[9]));
OAI21_X1 slo__sro_c374 (.ZN (n_10), .A (slo__sro_n552), .B1 (slo__sro_n553), .B2 (slo__sro_n551));
XNOR2_X1 slo__sro_c375 (.ZN (slo__sro_n550), .A (p_0[9]), .B (Multiplier[9]));
XNOR2_X1 slo__sro_c376 (.ZN (p_1[9]), .A (slo__sro_n550), .B (CLOCK_slo__sro_n1251));
XNOR2_X1 slo__sro_c507 (.ZN (p_1[11]), .A (slo__sro_n739), .B (n_11));
XNOR2_X1 slo__mro_c532 (.ZN (p_1[19]), .A (slo__mro_n781), .B (n_19));
INV_X1 slo__xsl_c482 (.ZN (slo__xsl_n703), .A (slo__sro_n326));
INV_X1 slo__xsl_c483 (.ZN (slo__xsl_n702), .A (slo__xsl_n703));
XNOR2_X1 slo__mro_c490 (.ZN (p_1[12]), .A (slo__sro_n57), .B (n_12));
NAND2_X1 slo__sro_c503 (.ZN (slo__sro_n741), .A1 (p_0[11]), .A2 (Multiplier[11]));
NOR2_X1 slo__sro_c504 (.ZN (slo__sro_n740), .A1 (p_0[11]), .A2 (Multiplier[11]));
OAI21_X1 slo__sro_c505 (.ZN (n_12), .A (slo__sro_n741), .B1 (slo__sro_n742), .B2 (slo__sro_n740));
NOR2_X1 slo__sro_c551 (.ZN (slo__sro_n814), .A1 (slo__sro_n186), .A2 (Multiplier[27]));
OAI21_X1 slo__sro_c552 (.ZN (n_28), .A (slo__sro_n815), .B1 (slo__sro_n814), .B2 (slo__sro_n816));
XNOR2_X2 slo__sro_c553 (.ZN (slo__sro_n813), .A (p_0[27]), .B (Multiplier[27]));
XNOR2_X1 slo__sro_c554 (.ZN (p_1[27]), .A (slo__sro_n813), .B (slo__sro_n186));
XNOR2_X1 slo__mro_c597 (.ZN (p_1[15]), .A (slo__mro_n862), .B (n_15));
NOR2_X1 slo__mro_c579 (.ZN (slo__sro_n101), .A1 (p_0[14]), .A2 (Multiplier[14]));
OAI21_X1 slo__sro_c609 (.ZN (n_19), .A (slo__sro_n879), .B1 (slo__sro_n880), .B2 (slo__sro_n878));
XNOR2_X2 slo__sro_c610 (.ZN (slo__sro_n877), .A (p_0[18]), .B (Multiplier[18]));
XNOR2_X2 slo__sro_c611 (.ZN (p_1[18]), .A (slo__sro_n877), .B (slo__sro_n157));
XNOR2_X2 CLOCK_slo__mro_c736 (.ZN (p_1[4]), .A (CLOCK_slo__mro_n1145), .B (n_4));
NAND2_X1 CLOCK_slo__sro_c749 (.ZN (CLOCK_slo__sro_n1160), .A1 (CLOCK_slo__sro_n1161), .A2 (CLOCK_slo__sro_n1162));
OR2_X1 CLOCK_slo__sro_c750 (.ZN (CLOCK_slo__sro_n1159), .A1 (p_0[30]), .A2 (n_34));
OAI21_X1 CLOCK_slo__sro_c751 (.ZN (CLOCK_slo__sro_n1158), .A (CLOCK_slo__sro_n1160)
    , .B1 (n_32), .B2 (CLOCK_slo__sro_n1159));
NAND2_X1 CLOCK_slo__sro_c788 (.ZN (CLOCK_slo__sro_n1194), .A1 (p_0[22]), .A2 (Multiplier[22]));
NOR2_X2 CLOCK_slo__mro_c781 (.ZN (CLOCK_slo__mro_n1184), .A1 (p_0[3]), .A2 (Multiplier[3]));
OAI21_X1 CLOCK_slo__sro_c790 (.ZN (n_23), .A (CLOCK_slo__sro_n1194), .B1 (CLOCK_slo__sro_n1195), .B2 (CLOCK_slo__sro_n1193));
XNOR2_X2 CLOCK_slo__sro_c791 (.ZN (CLOCK_slo__sro_n1192), .A (p_0[22]), .B (Multiplier[22]));
XNOR2_X2 CLOCK_slo__sro_c792 (.ZN (p_1[22]), .A (CLOCK_slo__sro_n1192), .B (CLOCK_slo__sro_n1270));
OAI21_X1 CLOCK_slo__sro_c814 (.ZN (CLOCK_slo__sro_n1225), .A (n_28), .B1 (p_0[28]), .B2 (Multiplier[28]));
NAND2_X1 CLOCK_slo__sro_c815 (.ZN (CLOCK_slo__sro_n1224), .A1 (CLOCK_slo__sro_n1225), .A2 (CLOCK_slo__sro_n1226));
XNOR2_X1 CLOCK_slo__sro_c816 (.ZN (CLOCK_slo__sro_n1223), .A (n_28), .B (Multiplier[28]));
XNOR2_X1 CLOCK_slo__sro_c817 (.ZN (p_1[28]), .A (CLOCK_slo__sro_n1223), .B (p_0[28]));
NAND2_X1 CLOCK_slo__sro_c839 (.ZN (CLOCK_slo__sro_n1253), .A1 (p_0[8]), .A2 (Multiplier[8]));
NOR2_X1 CLOCK_slo__sro_c840 (.ZN (CLOCK_slo__sro_n1252), .A1 (p_0[8]), .A2 (Multiplier[8]));
OAI21_X1 CLOCK_slo__sro_c841 (.ZN (CLOCK_slo__sro_n1251), .A (CLOCK_slo__sro_n1253)
    , .B1 (CLOCK_slo__sro_n1254), .B2 (CLOCK_slo__sro_n1252));
XNOR2_X1 CLOCK_slo__sro_c842 (.ZN (CLOCK_slo__sro_n1250), .A (p_0[8]), .B (Multiplier[8]));
XNOR2_X1 CLOCK_slo__sro_c843 (.ZN (p_1[8]), .A (CLOCK_slo__sro_n1250), .B (n_8));
OAI21_X1 CLOCK_slo__sro_c855 (.ZN (CLOCK_slo__sro_n1271), .A (slo__sro_n142), .B1 (p_0[21]), .B2 (Multiplier[21]));
NAND2_X1 CLOCK_slo__sro_c856 (.ZN (CLOCK_slo__sro_n1270), .A1 (CLOCK_slo__sro_n1271), .A2 (CLOCK_slo__sro_n1272));
XNOR2_X1 CLOCK_slo__sro_c857 (.ZN (CLOCK_slo__sro_n1269), .A (p_0[21]), .B (Multiplier[21]));
XNOR2_X1 CLOCK_slo__sro_c858 (.ZN (p_1[21]), .A (CLOCK_slo__sro_n1269), .B (slo__sro_n142));
OAI22_X1 CLOCK_slo__sro_c876 (.ZN (CLOCK_slo__sro_n1294), .A1 (n_33), .A2 (Multiplier[30])
    , .B1 (p_0[30]), .B2 (n_34));
NAND2_X1 CLOCK_slo__sro_c929 (.ZN (CLOCK_slo__sro_n1409), .A1 (n_2), .A2 (p_0[2]));
NAND3_X1 CLOCK_slo__sro_c930 (.ZN (n_3), .A1 (CLOCK_slo__sro_n1409), .A2 (CLOCK_slo__sro_n1410), .A3 (CLOCK_slo__sro_n1411));
XNOR2_X1 CLOCK_slo__sro_c931 (.ZN (CLOCK_slo__sro_n1408), .A (p_0[2]), .B (Multiplier[2]));
XNOR2_X1 CLOCK_slo__sro_c932 (.ZN (p_1[2]), .A (CLOCK_slo__sro_n1408), .B (n_2));

endmodule //datapath__0_191

module datapath__0_187 (opt_ipoPP_1, p_0, p_1, p_2);

output [31:0] p_2;
input [31:0] p_0;
input [31:0] p_1;
input opt_ipoPP_1;
wire slo__sro_n845;
wire slo__sro_n516;
wire n_1;
wire n_2;
wire n_4;
wire n_5;
wire n_6;
wire n_8;
wire n_9;
wire n_10;
wire n_12;
wire n_13;
wire n_14;
wire n_15;
wire n_16;
wire n_17;
wire n_19;
wire n_20;
wire n_21;
wire n_24;
wire n_25;
wire n_27;
wire n_28;
wire n_29;
wire n_30;
wire n_32;
wire n_0;
wire n_34;
wire slo__sro_n160;
wire slo__sro_n161;
wire slo__sro_n162;
wire slo__sro_n163;
wire slo__sro_n164;
wire slo__sro_n202;
wire slo__sro_n203;
wire slo__sro_n204;
wire slo__sro_n205;
wire slo__sro_n92;
wire slo__sro_n93;
wire slo__sro_n94;
wire slo__sro_n95;
wire slo__sro_n130;
wire slo__sro_n131;
wire slo__sro_n132;
wire slo__sro_n133;
wire slo__sro_n134;
wire slo__sro_n259;
wire slo__sro_n260;
wire slo__sro_n261;
wire slo__sro_n262;
wire slo__sro_n289;
wire slo__sro_n290;
wire slo__sro_n291;
wire slo__sro_n292;
wire slo__sro_n448;
wire slo__sro_n449;
wire slo__sro_n450;
wire slo__sro_n451;
wire slo__sro_n452;
wire slo__sro_n517;
wire slo__sro_n518;
wire slo__sro_n519;
wire slo__sro_n568;
wire slo__sro_n569;
wire slo__sro_n570;
wire slo__sro_n571;
wire slo__sro_n572;
wire slo__sro_n731;
wire slo__sro_n732;
wire slo__sro_n733;
wire slo__sro_n734;
wire slo__sro_n735;
wire slo__sro_n846;
wire slo__sro_n847;
wire slo__sro_n848;
wire slo__sro_n849;
wire CLOCK_slo__sro_n1046;
wire CLOCK_slo__sro_n1047;
wire CLOCK_slo__sro_n1048;
wire CLOCK_slo__sro_n1049;
wire CLOCK_slo__sro_n1080;
wire CLOCK_slo__sro_n1081;
wire CLOCK_slo__sro_n1082;
wire CLOCK_slo__sro_n1083;
wire CLOCK_slo__sro_n1084;
wire CLOCK_slo__sro_n1109;
wire CLOCK_slo__sro_n1110;
wire CLOCK_slo__sro_n1111;
wire CLOCK_slo__sro_n1112;
wire CLOCK_slo__sro_n1113;
wire CLOCK_slo__sro_n1156;


INV_X1 i_36 (.ZN (n_34), .A (p_0[30]));
INV_X2 i_34 (.ZN (n_32), .A (n_30));
XNOR2_X1 CLOCK_slo__sro_c1164 (.ZN (p_2[30]), .A (n_32), .B (n_0));
OAI22_X1 i_31 (.ZN (n_0), .A1 (n_34), .A2 (opt_ipoPP_1), .B1 (p_0[30]), .B2 (p_1[30]));
FA_X1 i_30 (.CO (n_30), .S (p_2[29]), .A (p_0[29]), .B (p_1[29]), .CI (n_29));
FA_X1 i_29 (.CO (n_29), .S (p_2[28]), .A (p_0[28]), .B (p_1[28]), .CI (n_28));
FA_X1 i_28 (.CO (n_28), .S (p_2[27]), .A (p_0[27]), .B (p_1[27]), .CI (n_27));
FA_X1 i_27 (.CO (n_27), .S (p_2[26]), .A (p_0[26]), .B (p_1[26]), .CI (slo__sro_n569));
INV_X1 slo__sro_c500 (.ZN (slo__sro_n735), .A (p_1[10]));
FA_X1 i_25 (.CO (n_25), .S (p_2[24]), .A (p_0[24]), .B (p_1[24]), .CI (n_24));
FA_X1 i_24 (.CO (n_24), .S (p_2[23]), .A (p_0[23]), .B (p_1[23]), .CI (slo__sro_n131));
NOR2_X1 slo__sro_c193 (.ZN (slo__sro_n260), .A1 (p_1[9]), .A2 (p_0[9]));
INV_X1 CLOCK_slo__sro_c776 (.ZN (CLOCK_slo__sro_n1113), .A (n_2));
FA_X1 i_21 (.CO (n_21), .S (p_2[20]), .A (p_0[20]), .B (p_1[20]), .CI (n_20));
FA_X1 i_20 (.CO (n_20), .S (p_2[19]), .A (p_0[19]), .B (p_1[19]), .CI (n_19));
INV_X1 slo__sro_c191 (.ZN (slo__sro_n262), .A (n_9));
INV_X1 slo__sro_c136 (.ZN (slo__sro_n205), .A (slo__sro_n161));
INV_X1 CLOCK_slo__sro_c749 (.ZN (CLOCK_slo__sro_n1084), .A (n_21));
FA_X1 i_16 (.CO (n_16), .S (p_2[15]), .A (p_0[15]), .B (p_1[15]), .CI (n_15));
FA_X1 i_15 (.CO (n_15), .S (p_2[14]), .A (p_0[14]), .B (p_1[14]), .CI (n_14));
NOR2_X1 slo__sro_c410 (.ZN (slo__sro_n570), .A1 (p_1[25]), .A2 (p_0[25]));
INV_X2 slo__sro_c69 (.ZN (slo__sro_n134), .A (CLOCK_slo__sro_n1081));
FA_X1 i_12 (.CO (n_12), .S (p_2[11]), .A (p_0[11]), .B (p_1[11]), .CI (slo__sro_n732));
INV_X1 slo__sro_c575 (.ZN (slo__sro_n849), .A (n_30));
INV_X1 slo__sro_c220 (.ZN (slo__sro_n292), .A (slo__sro_n449));
FA_X1 i_9 (.CO (n_9), .S (p_2[8]), .A (p_0[8]), .B (p_1[8]), .CI (n_8));
INV_X1 slo__sro_c375 (.ZN (slo__sro_n519), .A (n_13));
NAND2_X1 slo__sro_c376 (.ZN (slo__sro_n518), .A1 (p_1[13]), .A2 (p_0[13]));
FA_X1 i_6 (.CO (n_6), .S (p_2[5]), .A (p_0[5]), .B (p_1[5]), .CI (n_5));
FA_X1 i_5 (.CO (n_5), .S (p_2[4]), .A (p_0[4]), .B (p_1[4]), .CI (n_4));
FA_X1 i_4 (.CO (n_4), .S (p_2[3]), .A (p_0[3]), .B (p_1[3]), .CI (CLOCK_slo__sro_n1110));
FA_X1 i_2 (.CO (n_2), .S (p_2[1]), .A (p_0[1]), .B (p_1[1]), .CI (n_1));
HA_X1 i_1 (.CO (n_1), .S (p_2[0]), .A (p_0[0]), .B (p_1[0]));
INV_X1 slo__sro_c96 (.ZN (slo__sro_n164), .A (n_17));
NAND2_X1 slo__sro_c97 (.ZN (slo__sro_n163), .A1 (p_1[17]), .A2 (p_0[17]));
NOR2_X1 slo__sro_c98 (.ZN (slo__sro_n162), .A1 (p_1[17]), .A2 (p_0[17]));
OAI21_X1 slo__sro_c99 (.ZN (slo__sro_n161), .A (slo__sro_n163), .B1 (slo__sro_n164), .B2 (slo__sro_n162));
XNOR2_X1 slo__sro_c100 (.ZN (slo__sro_n160), .A (p_1[17]), .B (p_0[17]));
XNOR2_X1 slo__sro_c101 (.ZN (p_2[17]), .A (n_17), .B (slo__sro_n160));
NAND2_X1 slo__sro_c137 (.ZN (slo__sro_n204), .A1 (p_1[18]), .A2 (p_0[18]));
NOR2_X1 slo__sro_c138 (.ZN (slo__sro_n203), .A1 (p_1[18]), .A2 (p_0[18]));
OAI21_X1 slo__sro_c139 (.ZN (n_19), .A (slo__sro_n204), .B1 (slo__sro_n205), .B2 (slo__sro_n203));
XNOR2_X1 slo__sro_c140 (.ZN (slo__sro_n202), .A (p_1[18]), .B (p_0[18]));
XNOR2_X1 slo__sro_c141 (.ZN (p_2[18]), .A (slo__sro_n202), .B (slo__sro_n161));
NAND2_X1 slo__sro_c192 (.ZN (slo__sro_n261), .A1 (p_1[9]), .A2 (p_0[9]));
INV_X1 slo__sro_c29 (.ZN (slo__sro_n95), .A (n_12));
NAND2_X1 slo__sro_c30 (.ZN (slo__sro_n94), .A1 (p_1[12]), .A2 (p_0[12]));
NOR2_X1 slo__sro_c31 (.ZN (slo__sro_n93), .A1 (p_1[12]), .A2 (p_0[12]));
OAI21_X2 slo__sro_c32 (.ZN (n_13), .A (slo__sro_n94), .B1 (slo__sro_n95), .B2 (slo__sro_n93));
XNOR2_X1 slo__sro_c33 (.ZN (slo__sro_n92), .A (p_1[12]), .B (p_0[12]));
XNOR2_X1 slo__sro_c34 (.ZN (p_2[12]), .A (n_12), .B (slo__sro_n92));
NAND2_X1 slo__sro_c70 (.ZN (slo__sro_n133), .A1 (p_1[22]), .A2 (p_0[22]));
NOR2_X1 slo__sro_c71 (.ZN (slo__sro_n132), .A1 (p_1[22]), .A2 (p_0[22]));
OAI21_X1 slo__sro_c72 (.ZN (slo__sro_n131), .A (slo__sro_n133), .B1 (slo__sro_n134), .B2 (slo__sro_n132));
XNOR2_X1 slo__sro_c73 (.ZN (slo__sro_n130), .A (p_1[22]), .B (p_0[22]));
XNOR2_X1 slo__sro_c74 (.ZN (p_2[22]), .A (slo__sro_n130), .B (CLOCK_slo__sro_n1081));
OAI21_X2 slo__sro_c194 (.ZN (n_10), .A (slo__sro_n261), .B1 (slo__sro_n260), .B2 (slo__sro_n262));
XNOR2_X1 slo__sro_c195 (.ZN (slo__sro_n259), .A (p_1[9]), .B (p_0[9]));
XNOR2_X1 slo__sro_c196 (.ZN (p_2[9]), .A (slo__sro_n259), .B (n_9));
NAND2_X1 slo__sro_c221 (.ZN (slo__sro_n291), .A1 (p_1[7]), .A2 (p_0[7]));
NOR2_X1 slo__sro_c222 (.ZN (slo__sro_n290), .A1 (p_1[7]), .A2 (p_0[7]));
OAI21_X1 slo__sro_c223 (.ZN (n_8), .A (slo__sro_n291), .B1 (slo__sro_n292), .B2 (slo__sro_n290));
XNOR2_X1 slo__sro_c224 (.ZN (slo__sro_n289), .A (p_1[7]), .B (p_0[7]));
XNOR2_X1 slo__sro_c225 (.ZN (p_2[7]), .A (slo__sro_n449), .B (slo__sro_n289));
INV_X1 slo__sro_c319 (.ZN (slo__sro_n452), .A (n_6));
NAND2_X1 slo__sro_c320 (.ZN (slo__sro_n451), .A1 (p_1[6]), .A2 (p_0[6]));
NOR2_X1 slo__sro_c321 (.ZN (slo__sro_n450), .A1 (p_1[6]), .A2 (p_0[6]));
OAI21_X1 slo__sro_c322 (.ZN (slo__sro_n449), .A (slo__sro_n451), .B1 (slo__sro_n452), .B2 (slo__sro_n450));
XNOR2_X1 slo__sro_c323 (.ZN (slo__sro_n448), .A (p_1[6]), .B (p_0[6]));
XNOR2_X1 slo__sro_c324 (.ZN (p_2[6]), .A (n_6), .B (slo__sro_n448));
NOR2_X1 slo__sro_c377 (.ZN (slo__sro_n517), .A1 (p_1[13]), .A2 (p_0[13]));
OAI21_X1 slo__sro_c378 (.ZN (n_14), .A (slo__sro_n518), .B1 (slo__sro_n519), .B2 (slo__sro_n517));
XNOR2_X1 slo__sro_c379 (.ZN (slo__sro_n516), .A (p_1[13]), .B (p_0[13]));
XNOR2_X1 slo__sro_c380 (.ZN (p_2[13]), .A (slo__sro_n516), .B (n_13));
INV_X2 slo__sro_c408 (.ZN (slo__sro_n572), .A (n_25));
NAND2_X1 slo__sro_c409 (.ZN (slo__sro_n571), .A1 (p_1[25]), .A2 (p_0[25]));
OAI21_X2 slo__sro_c411 (.ZN (slo__sro_n569), .A (slo__sro_n571), .B1 (slo__sro_n572), .B2 (slo__sro_n570));
XNOR2_X1 slo__sro_c412 (.ZN (slo__sro_n568), .A (p_1[25]), .B (p_0[25]));
XNOR2_X1 slo__sro_c413 (.ZN (p_2[25]), .A (n_25), .B (slo__sro_n568));
NAND2_X1 slo__sro_c501 (.ZN (slo__sro_n734), .A1 (n_10), .A2 (p_0[10]));
NOR2_X2 slo__sro_c502 (.ZN (slo__sro_n733), .A1 (n_10), .A2 (p_0[10]));
OAI21_X1 slo__sro_c503 (.ZN (slo__sro_n732), .A (slo__sro_n734), .B1 (slo__sro_n733), .B2 (slo__sro_n735));
XNOR2_X2 slo__sro_c504 (.ZN (slo__sro_n731), .A (p_1[10]), .B (p_0[10]));
XNOR2_X1 slo__sro_c505 (.ZN (p_2[10]), .A (slo__sro_n731), .B (n_10));
NOR2_X1 slo__sro_c576 (.ZN (slo__sro_n848), .A1 (p_1[30]), .A2 (p_0[30]));
NAND2_X1 slo__sro_c577 (.ZN (slo__sro_n847), .A1 (slo__sro_n848), .A2 (slo__sro_n849));
OR2_X1 slo__sro_c578 (.ZN (slo__sro_n846), .A1 (opt_ipoPP_1), .A2 (n_34));
OAI21_X1 slo__sro_c579 (.ZN (slo__sro_n845), .A (slo__sro_n847), .B1 (n_32), .B2 (slo__sro_n846));
INV_X1 CLOCK_slo__sro_c713 (.ZN (CLOCK_slo__sro_n1049), .A (n_16));
NAND2_X1 CLOCK_slo__sro_c714 (.ZN (CLOCK_slo__sro_n1048), .A1 (p_1[16]), .A2 (p_0[16]));
NOR2_X1 CLOCK_slo__sro_c715 (.ZN (CLOCK_slo__sro_n1047), .A1 (p_1[16]), .A2 (p_0[16]));
OAI21_X1 CLOCK_slo__sro_c716 (.ZN (n_17), .A (CLOCK_slo__sro_n1048), .B1 (CLOCK_slo__sro_n1049), .B2 (CLOCK_slo__sro_n1047));
XNOR2_X1 CLOCK_slo__sro_c717 (.ZN (CLOCK_slo__sro_n1046), .A (p_1[16]), .B (p_0[16]));
XNOR2_X1 CLOCK_slo__sro_c718 (.ZN (p_2[16]), .A (CLOCK_slo__sro_n1046), .B (n_16));
NAND2_X1 CLOCK_slo__sro_c750 (.ZN (CLOCK_slo__sro_n1083), .A1 (p_1[21]), .A2 (p_0[21]));
NOR2_X1 CLOCK_slo__sro_c751 (.ZN (CLOCK_slo__sro_n1082), .A1 (p_1[21]), .A2 (p_0[21]));
OAI21_X2 CLOCK_slo__sro_c752 (.ZN (CLOCK_slo__sro_n1081), .A (CLOCK_slo__sro_n1083)
    , .B1 (CLOCK_slo__sro_n1084), .B2 (CLOCK_slo__sro_n1082));
XNOR2_X1 CLOCK_slo__sro_c753 (.ZN (CLOCK_slo__sro_n1080), .A (p_1[21]), .B (p_0[21]));
XNOR2_X1 CLOCK_slo__sro_c754 (.ZN (p_2[21]), .A (CLOCK_slo__sro_n1080), .B (n_21));
NAND2_X1 CLOCK_slo__sro_c777 (.ZN (CLOCK_slo__sro_n1112), .A1 (p_1[2]), .A2 (p_0[2]));
NOR2_X1 CLOCK_slo__sro_c778 (.ZN (CLOCK_slo__sro_n1111), .A1 (p_1[2]), .A2 (p_0[2]));
OAI21_X1 CLOCK_slo__sro_c779 (.ZN (CLOCK_slo__sro_n1110), .A (CLOCK_slo__sro_n1112)
    , .B1 (CLOCK_slo__sro_n1111), .B2 (CLOCK_slo__sro_n1113));
XNOR2_X1 CLOCK_slo__sro_c780 (.ZN (CLOCK_slo__sro_n1109), .A (p_1[2]), .B (p_0[2]));
XNOR2_X1 CLOCK_slo__sro_c781 (.ZN (p_2[2]), .A (CLOCK_slo__sro_n1109), .B (n_2));
INV_X1 CLOCK_slo__sro_c824 (.ZN (CLOCK_slo__sro_n1156), .A (p_0[31]));
XNOR2_X1 CLOCK_slo__sro_c825 (.ZN (p_2[31]), .A (slo__sro_n845), .B (CLOCK_slo__sro_n1156));

endmodule //datapath__0_187

module datapath__0_186 (p_0_8_PP_0, opt_ipoPP_0, opt_ipoPP_2, Multiplier, p_0, p_1);

output [31:0] p_1;
input [31:0] Multiplier;
input [31:0] p_0;
input p_0_8_PP_0;
input opt_ipoPP_0;
input opt_ipoPP_2;
wire slo_n811;
wire slo__sro_n608;
wire n_1;
wire n_2;
wire n_3;
wire n_4;
wire n_5;
wire n_6;
wire n_8;
wire n_10;
wire n_11;
wire n_13;
wire CLOCK_slo__sro_n1518;
wire n_15;
wire n_16;
wire n_18;
wire n_19;
wire n_20;
wire n_22;
wire n_25;
wire n_26;
wire n_28;
wire n_29;
wire n_30;
wire n_32;
wire n_0;
wire n_34;
wire CLOCK_slo__sro_n1460;
wire n_31;
wire slo__sro_n57;
wire slo__sro_n58;
wire slo__sro_n59;
wire slo__sro_n60;
wire slo__sro_n98;
wire slo__sro_n99;
wire slo__sro_n100;
wire slo__sro_n101;
wire slo__sro_n111;
wire slo__sro_n112;
wire slo__sro_n113;
wire slo__sro_n114;
wire slo__sro_n115;
wire slo__sro_n140;
wire slo__sro_n141;
wire slo__sro_n142;
wire slo__sro_n143;
wire slo__sro_n144;
wire slo__sro_n157;
wire slo__sro_n158;
wire slo__sro_n159;
wire slo__sro_n160;
wire slo__sro_n172;
wire slo__sro_n173;
wire slo__sro_n174;
wire slo__sro_n175;
wire slo__sro_n176;
wire CLOCK_slo__sro_n1517;
wire slo__sro_n190;
wire slo__sro_n191;
wire slo__sro_n192;
wire slo__sro_n193;
wire slo__sro_n210;
wire slo__sro_n211;
wire slo__sro_n212;
wire slo__sro_n213;
wire slo__sro_n241;
wire slo__sro_n242;
wire slo__sro_n243;
wire slo__sro_n244;
wire slo__sro_n245;
wire slo__sro_n409;
wire slo__sro_n410;
wire slo__sro_n411;
wire slo__sro_n412;
wire slo__sro_n424;
wire slo__sro_n425;
wire slo__sro_n426;
wire slo__sro_n427;
wire slo__sro_n475;
wire slo__sro_n476;
wire slo__sro_n477;
wire slo__sro_n478;
wire slo__sro_n609;
wire slo__sro_n610;
wire slo__sro_n611;
wire slo__sro_n504;
wire slo__sro_n505;
wire slo__sro_n506;
wire slo__sro_n507;
wire slo__sro_n508;
wire slo__sro_n623;
wire slo__sro_n624;
wire slo__sro_n625;
wire slo__sro_n626;
wire slo__sro_n815;
wire slo__sro_n816;
wire slo__sro_n817;
wire slo__sro_n818;
wire slo__sro_n819;
wire slo__sro_n832;
wire slo__sro_n833;
wire slo__sro_n834;
wire slo__sro_n835;
wire slo__sro_n900;
wire slo__sro_n901;
wire slo__sro_n902;
wire slo__sro_n903;
wire slo__mro_n915;
wire CLOCK_slo__sro_n1461;
wire CLOCK_slo__sro_n1462;
wire CLOCK_slo__sro_n1463;
wire CLOCK_slo__mro_n1443;
wire CLOCK_slo__mro_n1444;
wire CLOCK_slo__sro_n1519;
wire CLOCK_slo__sro_n1783;
wire CLOCK_slo__sro_n1784;
wire CLOCK_slo__sro_n1785;


INV_X1 i_36 (.ZN (n_34), .A (Multiplier[30]));
NAND2_X1 CLOCK_slo__sro_c1144 (.ZN (CLOCK_slo__sro_n1519), .A1 (slo__sro_n242), .A2 (Multiplier[27]));
INV_X1 i_34 (.ZN (n_32), .A (n_30));
OAI33_X1 i_33 (.ZN (n_31), .A1 (n_32), .A2 (opt_ipoPP_2), .A3 (n_34), .B1 (n_30), .B2 (p_0[30]), .B3 (Multiplier[30]));
XOR2_X1 i_32 (.Z (p_1[31]), .A (Multiplier[31]), .B (n_31));
OAI22_X1 i_31 (.ZN (n_0), .A1 (n_34), .A2 (opt_ipoPP_2), .B1 (Multiplier[30]), .B2 (p_0[30]));
XNOR2_X1 i_0 (.ZN (p_1[30]), .A (n_32), .B (n_0));
FA_X1 i_30 (.CO (n_30), .S (p_1[29]), .A (Multiplier[29]), .B (p_0[29]), .CI (n_29));
INV_X1 slo__sro_c681 (.ZN (slo__sro_n903), .A (p_0[10]));
INV_X1 slo__sro_c472 (.ZN (slo__sro_n611), .A (p_0[9]));
NAND2_X1 slo__sro_c619 (.ZN (slo__sro_n818), .A1 (p_0[23]), .A2 (Multiplier[23]));
FA_X1 i_25 (.CO (n_25), .S (p_1[24]), .A (Multiplier[24]), .B (p_0[24]), .CI (slo__sro_n816));
INV_X1 slo__sro_c632 (.ZN (slo__sro_n835), .A (n_28));
INV_X1 slo__sro_c96 (.ZN (slo__sro_n160), .A (n_4));
OAI21_X1 CLOCK_slo__sro_c1145 (.ZN (CLOCK_slo__sro_n1518), .A (p_0[27]), .B1 (slo__sro_n242), .B2 (Multiplier[27]));
INV_X1 slo__sro_c168 (.ZN (slo__sro_n245), .A (n_26));
INV_X1 slo__sro_c55 (.ZN (slo__sro_n115), .A (n_6));
FA_X1 i_19 (.CO (n_19), .S (p_1[18]), .A (Multiplier[18]), .B (p_0[18]), .CI (n_18));
FA_X1 i_18 (.CO (n_18), .S (p_1[17]), .A (Multiplier[17]), .B (p_0[17]), .CI (slo__sro_n173));
NAND2_X1 slo__sro_c124 (.ZN (slo__sro_n193), .A1 (p_0[13]), .A2 (Multiplier[13]));
FA_X1 i_16 (.CO (n_16), .S (p_1[15]), .A (Multiplier[15]), .B (p_0[15]), .CI (n_15));
FA_X1 i_15 (.CO (n_15), .S (p_1[14]), .A (Multiplier[14]), .B (p_0[14]), .CI (slo__sro_n190));
NAND2_X1 slo__sro_c141 (.ZN (slo__sro_n213), .A1 (p_0[20]), .A2 (Multiplier[20]));
INV_X2 slo__sro_c41 (.ZN (slo__sro_n101), .A (n_19));
NAND2_X1 slo__sro_c489 (.ZN (slo__sro_n625), .A1 (p_0[25]), .A2 (Multiplier[25]));
XNOR2_X1 slo__mro_c695 (.ZN (slo__mro_n915), .A (n_13), .B (Multiplier[13]));
INV_X1 slo__sro_c488 (.ZN (slo__sro_n626), .A (n_25));
NAND2_X1 slo__sro_c473 (.ZN (slo__sro_n610), .A1 (slo__sro_n476), .A2 (Multiplier[9]));
INV_X1 slo__sro_c618 (.ZN (slo__sro_n819), .A (slo__sro_n141));
INV_X1 slo__sro_c82 (.ZN (slo__sro_n144), .A (n_22));
INV_X1 slo__sro_c110 (.ZN (slo__sro_n176), .A (n_16));
NAND2_X1 slo__sro_c315 (.ZN (slo__sro_n426), .A1 (slo__sro_n112), .A2 (Multiplier[7]));
FA_X1 i_3 (.CO (n_3), .S (p_1[2]), .A (Multiplier[2]), .B (p_0[2]), .CI (n_2));
FA_X1 i_2 (.CO (n_2), .S (p_1[1]), .A (Multiplier[1]), .B (p_0[1]), .CI (n_1));
HA_X1 i_1 (.CO (n_1), .S (p_1[0]), .A (Multiplier[0]), .B (p_0[0]));
INV_X1 slo__sro_c1 (.ZN (slo__sro_n60), .A (slo__sro_n505));
NAND2_X1 slo__sro_c2 (.ZN (slo__sro_n59), .A1 (p_0[12]), .A2 (Multiplier[12]));
NOR2_X1 slo__sro_c3 (.ZN (slo__sro_n58), .A1 (p_0[12]), .A2 (Multiplier[12]));
OAI21_X2 slo__sro_c4 (.ZN (n_13), .A (slo__sro_n59), .B1 (slo__sro_n58), .B2 (slo__sro_n60));
XNOR2_X2 slo__sro_c5 (.ZN (slo__sro_n57), .A (p_0[12]), .B (Multiplier[12]));
XNOR2_X1 slo__sro_c6 (.ZN (p_1[12]), .A (slo__sro_n57), .B (slo__sro_n505));
NAND2_X1 slo__sro_c42 (.ZN (slo__sro_n100), .A1 (p_0[19]), .A2 (Multiplier[19]));
NOR2_X1 slo__sro_c43 (.ZN (slo__sro_n99), .A1 (p_0[19]), .A2 (Multiplier[19]));
OAI21_X1 slo__sro_c44 (.ZN (n_20), .A (slo__sro_n100), .B1 (slo__sro_n101), .B2 (slo__sro_n99));
XNOR2_X1 slo__sro_c45 (.ZN (slo__sro_n98), .A (p_0[19]), .B (Multiplier[19]));
XNOR2_X1 slo__sro_c46 (.ZN (p_1[19]), .A (n_19), .B (slo__sro_n98));
NAND2_X1 slo__sro_c56 (.ZN (slo__sro_n114), .A1 (p_0[6]), .A2 (Multiplier[6]));
NOR2_X2 slo__sro_c57 (.ZN (slo__sro_n113), .A1 (p_0[6]), .A2 (Multiplier[6]));
OAI21_X2 slo__sro_c58 (.ZN (slo__sro_n112), .A (slo__sro_n114), .B1 (slo__sro_n115), .B2 (slo__sro_n113));
XNOR2_X1 slo__sro_c59 (.ZN (slo__sro_n111), .A (p_0[6]), .B (Multiplier[6]));
XNOR2_X1 slo__sro_c60 (.ZN (p_1[6]), .A (slo__sro_n111), .B (n_6));
NAND2_X1 slo__sro_c83 (.ZN (slo__sro_n143), .A1 (p_0[22]), .A2 (Multiplier[22]));
NOR2_X1 slo__sro_c84 (.ZN (slo__sro_n142), .A1 (p_0[22]), .A2 (Multiplier[22]));
OAI21_X2 slo__sro_c85 (.ZN (slo__sro_n141), .A (slo__sro_n143), .B1 (slo__sro_n144), .B2 (slo__sro_n142));
XNOR2_X2 slo__sro_c86 (.ZN (slo__sro_n140), .A (p_0[22]), .B (Multiplier[22]));
XNOR2_X2 slo__sro_c87 (.ZN (p_1[22]), .A (slo__sro_n140), .B (n_22));
NAND2_X1 slo__sro_c97 (.ZN (slo__sro_n159), .A1 (p_0[4]), .A2 (Multiplier[4]));
NOR2_X1 slo__sro_c98 (.ZN (slo__sro_n158), .A1 (p_0[4]), .A2 (Multiplier[4]));
OAI21_X1 slo__sro_c99 (.ZN (n_5), .A (slo__sro_n159), .B1 (slo__sro_n158), .B2 (slo__sro_n160));
XNOR2_X2 slo__sro_c100 (.ZN (slo__sro_n157), .A (p_0[4]), .B (Multiplier[4]));
XNOR2_X2 slo__sro_c101 (.ZN (p_1[4]), .A (slo__sro_n157), .B (n_4));
NAND2_X1 slo__sro_c111 (.ZN (slo__sro_n175), .A1 (p_0[16]), .A2 (Multiplier[16]));
NOR2_X1 slo__sro_c112 (.ZN (slo__sro_n174), .A1 (p_0[16]), .A2 (Multiplier[16]));
OAI21_X1 slo__sro_c113 (.ZN (slo__sro_n173), .A (slo__sro_n175), .B1 (slo__sro_n176), .B2 (slo__sro_n174));
XNOR2_X1 slo__sro_c114 (.ZN (slo__sro_n172), .A (p_0[16]), .B (Multiplier[16]));
XNOR2_X1 slo__sro_c115 (.ZN (p_1[16]), .A (slo__sro_n172), .B (n_16));
NAND2_X1 slo__sro_c125 (.ZN (slo__sro_n192), .A1 (n_13), .A2 (Multiplier[13]));
NAND2_X1 slo__sro_c126 (.ZN (slo__sro_n191), .A1 (n_13), .A2 (p_0[13]));
NAND3_X1 slo__sro_c127 (.ZN (slo__sro_n190), .A1 (slo__sro_n192), .A2 (slo__sro_n191), .A3 (slo__sro_n193));
XNOR2_X1 CLOCK_slo__sro_c1092 (.ZN (p_1[21]), .A (CLOCK_slo__sro_n1460), .B (slo__sro_n210));
NAND2_X1 CLOCK_slo__sro_c1088 (.ZN (CLOCK_slo__sro_n1462), .A1 (p_0[21]), .A2 (Multiplier[21]));
NAND2_X1 slo__sro_c142 (.ZN (slo__sro_n212), .A1 (n_20), .A2 (Multiplier[20]));
NAND2_X1 slo__sro_c143 (.ZN (slo__sro_n211), .A1 (p_0[20]), .A2 (n_20));
NAND3_X1 slo__sro_c144 (.ZN (slo__sro_n210), .A1 (slo__sro_n213), .A2 (slo__sro_n211), .A3 (slo__sro_n212));
NAND2_X1 CLOCK_slo__sro_c1146 (.ZN (n_28), .A1 (CLOCK_slo__sro_n1518), .A2 (CLOCK_slo__sro_n1519));
XNOR2_X1 CLOCK_slo__sro_c1147 (.ZN (CLOCK_slo__sro_n1517), .A (slo__sro_n242), .B (Multiplier[27]));
NAND2_X1 slo__sro_c169 (.ZN (slo__sro_n244), .A1 (p_0[26]), .A2 (Multiplier[26]));
NOR2_X1 slo__sro_c170 (.ZN (slo__sro_n243), .A1 (p_0[26]), .A2 (Multiplier[26]));
OAI21_X1 slo__sro_c171 (.ZN (slo__sro_n242), .A (slo__sro_n244), .B1 (slo__sro_n245), .B2 (slo__sro_n243));
XNOR2_X2 slo__sro_c172 (.ZN (slo__sro_n241), .A (p_0[26]), .B (Multiplier[26]));
XNOR2_X2 slo__sro_c173 (.ZN (p_1[26]), .A (slo__sro_n241), .B (n_26));
NAND2_X1 slo__sro_c314 (.ZN (slo__sro_n427), .A1 (p_0[7]), .A2 (Multiplier[7]));
INV_X1 slo__sro_c298 (.ZN (slo__sro_n412), .A (n_3));
NAND2_X1 slo__sro_c299 (.ZN (slo__sro_n411), .A1 (p_0[3]), .A2 (Multiplier[3]));
NOR2_X1 slo__sro_c300 (.ZN (slo__sro_n410), .A1 (p_0[3]), .A2 (Multiplier[3]));
OAI21_X1 slo__sro_c301 (.ZN (n_4), .A (slo__sro_n411), .B1 (slo__sro_n410), .B2 (slo__sro_n412));
XNOR2_X2 slo__sro_c302 (.ZN (slo__sro_n409), .A (p_0[3]), .B (Multiplier[3]));
XNOR2_X2 slo__sro_c303 (.ZN (p_1[3]), .A (slo__sro_n409), .B (n_3));
NAND2_X1 slo__sro_c316 (.ZN (slo__sro_n425), .A1 (slo__sro_n112), .A2 (p_0[7]));
NAND3_X2 slo__sro_c317 (.ZN (n_8), .A1 (slo__sro_n425), .A2 (slo__sro_n426), .A3 (slo__sro_n427));
XNOR2_X2 slo__sro_c318 (.ZN (slo__sro_n424), .A (slo__sro_n112), .B (Multiplier[7]));
XNOR2_X2 slo__sro_c319 (.ZN (p_1[7]), .A (slo__sro_n424), .B (p_0[7]));
NAND2_X1 slo__sro_c351 (.ZN (slo__sro_n478), .A1 (n_8), .A2 (Multiplier[8]));
NOR2_X1 slo__sro_c352 (.ZN (slo__sro_n477), .A1 (n_8), .A2 (Multiplier[8]));
OAI21_X2 slo__sro_c353 (.ZN (slo__sro_n476), .A (slo__sro_n478), .B1 (slo_n811), .B2 (slo__sro_n477));
XNOR2_X1 slo__sro_c354 (.ZN (slo__sro_n475), .A (n_8), .B (Multiplier[8]));
XNOR2_X1 slo__sro_c355 (.ZN (p_1[8]), .A (slo__sro_n475), .B (p_0[8]));
NOR2_X1 slo__sro_c474 (.ZN (slo__sro_n609), .A1 (slo__sro_n476), .A2 (Multiplier[9]));
OAI21_X2 slo__sro_c475 (.ZN (n_10), .A (slo__sro_n610), .B1 (slo__sro_n609), .B2 (slo__sro_n611));
XNOR2_X1 slo__sro_c476 (.ZN (slo__sro_n608), .A (slo__sro_n476), .B (Multiplier[9]));
XNOR2_X1 slo__sro_c477 (.ZN (p_1[9]), .A (slo__sro_n608), .B (p_0[9]));
CLKBUF_X1 slo__L1_c1_c613 (.Z (slo_n811), .A (p_0_8_PP_0));
INV_X2 slo__sro_c380 (.ZN (slo__sro_n508), .A (n_11));
NAND2_X1 slo__sro_c381 (.ZN (slo__sro_n507), .A1 (p_0[11]), .A2 (Multiplier[11]));
NOR2_X2 slo__sro_c382 (.ZN (slo__sro_n506), .A1 (p_0[11]), .A2 (Multiplier[11]));
OAI21_X4 slo__sro_c383 (.ZN (slo__sro_n505), .A (slo__sro_n507), .B1 (slo__sro_n508), .B2 (slo__sro_n506));
XNOR2_X1 slo__sro_c384 (.ZN (slo__sro_n504), .A (p_0[11]), .B (Multiplier[11]));
XNOR2_X1 slo__sro_c385 (.ZN (p_1[11]), .A (n_11), .B (slo__sro_n504));
NOR2_X1 slo__sro_c490 (.ZN (slo__sro_n624), .A1 (p_0[25]), .A2 (Multiplier[25]));
OAI21_X1 slo__sro_c491 (.ZN (n_26), .A (slo__sro_n625), .B1 (slo__sro_n624), .B2 (slo__sro_n626));
XNOR2_X2 slo__sro_c492 (.ZN (slo__sro_n623), .A (p_0[25]), .B (Multiplier[25]));
XNOR2_X2 slo__sro_c493 (.ZN (p_1[25]), .A (slo__sro_n623), .B (n_25));
NOR2_X1 slo__sro_c620 (.ZN (slo__sro_n817), .A1 (p_0[23]), .A2 (Multiplier[23]));
OAI21_X1 slo__sro_c621 (.ZN (slo__sro_n816), .A (slo__sro_n818), .B1 (slo__sro_n817), .B2 (slo__sro_n819));
XNOR2_X1 slo__sro_c622 (.ZN (slo__sro_n815), .A (p_0[23]), .B (Multiplier[23]));
XNOR2_X2 slo__sro_c623 (.ZN (p_1[23]), .A (slo__sro_n815), .B (slo__sro_n141));
NAND2_X1 slo__sro_c633 (.ZN (slo__sro_n834), .A1 (p_0[28]), .A2 (Multiplier[28]));
NOR2_X1 slo__sro_c634 (.ZN (slo__sro_n833), .A1 (p_0[28]), .A2 (Multiplier[28]));
OAI21_X1 slo__sro_c635 (.ZN (n_29), .A (slo__sro_n834), .B1 (slo__sro_n833), .B2 (slo__sro_n835));
XNOR2_X1 slo__sro_c636 (.ZN (slo__sro_n832), .A (p_0[28]), .B (Multiplier[28]));
XNOR2_X1 slo__sro_c637 (.ZN (p_1[28]), .A (slo__sro_n832), .B (n_28));
NAND2_X1 slo__sro_c682 (.ZN (slo__sro_n902), .A1 (n_10), .A2 (Multiplier[10]));
NOR2_X1 slo__sro_c683 (.ZN (slo__sro_n901), .A1 (n_10), .A2 (Multiplier[10]));
OAI21_X2 slo__sro_c684 (.ZN (n_11), .A (slo__sro_n902), .B1 (slo__sro_n901), .B2 (slo__sro_n903));
XNOR2_X1 slo__sro_c685 (.ZN (slo__sro_n900), .A (n_10), .B (Multiplier[10]));
XNOR2_X1 slo__sro_c686 (.ZN (p_1[10]), .A (slo__sro_n900), .B (p_0[10]));
XNOR2_X1 slo__mro_c696 (.ZN (p_1[13]), .A (slo__mro_n915), .B (p_0[13]));
INV_X1 CLOCK_slo__sro_c1087 (.ZN (CLOCK_slo__sro_n1463), .A (slo__sro_n210));
NOR2_X1 CLOCK_slo__sro_c1089 (.ZN (CLOCK_slo__sro_n1461), .A1 (p_0[21]), .A2 (Multiplier[21]));
OAI21_X2 CLOCK_slo__sro_c1090 (.ZN (n_22), .A (CLOCK_slo__sro_n1462), .B1 (CLOCK_slo__sro_n1463), .B2 (CLOCK_slo__sro_n1461));
XNOR2_X1 CLOCK_slo__sro_c1091 (.ZN (CLOCK_slo__sro_n1460), .A (p_0[21]), .B (Multiplier[21]));
OAI21_X2 CLOCK_slo__mro_c1070 (.ZN (CLOCK_slo__mro_n1444), .A (slo__sro_n100), .B1 (slo__sro_n101), .B2 (slo__sro_n99));
XNOR2_X2 CLOCK_slo__mro_c1071 (.ZN (CLOCK_slo__mro_n1443), .A (CLOCK_slo__mro_n1444), .B (Multiplier[20]));
XNOR2_X1 CLOCK_slo__mro_c1072 (.ZN (p_1[20]), .A (CLOCK_slo__mro_n1443), .B (opt_ipoPP_0));
XNOR2_X1 CLOCK_slo__sro_c1148 (.ZN (p_1[27]), .A (CLOCK_slo__sro_n1517), .B (p_0[27]));
NAND2_X1 CLOCK_slo__sro_c1380 (.ZN (CLOCK_slo__sro_n1785), .A1 (p_0[5]), .A2 (Multiplier[5]));
OAI21_X1 CLOCK_slo__sro_c1381 (.ZN (CLOCK_slo__sro_n1784), .A (n_5), .B1 (p_0[5]), .B2 (Multiplier[5]));
NAND2_X2 CLOCK_slo__sro_c1382 (.ZN (n_6), .A1 (CLOCK_slo__sro_n1784), .A2 (CLOCK_slo__sro_n1785));
XNOR2_X1 CLOCK_slo__sro_c1383 (.ZN (CLOCK_slo__sro_n1783), .A (p_0[5]), .B (Multiplier[5]));
XNOR2_X1 CLOCK_slo__sro_c1384 (.ZN (p_1[5]), .A (CLOCK_slo__sro_n1783), .B (n_5));

endmodule //datapath__0_186

module datapath__0_182 (p_0, p_1, p_2);

output [31:0] p_2;
input [31:0] p_0;
input [31:0] p_1;
wire slo_n883;
wire CLOCK_slo__sro_n1336;
wire n_1;
wire n_2;
wire n_3;
wire n_4;
wire n_5;
wire n_6;
wire n_8;
wire n_9;
wire n_10;
wire n_11;
wire n_12;
wire n_13;
wire n_14;
wire n_16;
wire n_17;
wire n_18;
wire slo__sro_n756;
wire n_20;
wire n_21;
wire n_23;
wire slo__sro_n755;
wire n_25;
wire n_26;
wire n_27;
wire n_28;
wire n_30;
wire n_32;
wire n_0;
wire n_34;
wire n_33;
wire n_31;
wire slo__sro_n184;
wire slo__sro_n185;
wire slo__sro_n186;
wire slo__sro_n187;
wire slo__sro_n188;
wire slo__sro_n154;
wire slo__sro_n155;
wire slo__sro_n156;
wire slo__sro_n157;
wire slo__sro_n158;
wire slo__sro_n241;
wire slo__sro_n242;
wire slo__sro_n243;
wire slo__sro_n244;
wire slo__sro_n317;
wire slo__sro_n318;
wire slo__sro_n319;
wire slo__sro_n320;
wire slo__sro_n321;
wire slo__sro_n336;
wire slo__sro_n337;
wire slo__sro_n338;
wire slo__sro_n339;
wire slo__sro_n412;
wire slo__sro_n413;
wire slo__sro_n414;
wire slo__sro_n415;
wire slo__sro_n416;
wire slo__sro_n754;
wire slo__mro_n715;
wire slo__sro_n757;
wire slo__n898;
wire CLOCK_slo__sro_n1120;
wire CLOCK_slo__sro_n1121;
wire slo__sro_n503;
wire slo__sro_n504;
wire slo__sro_n505;
wire slo__sro_n506;
wire CLOCK_slo__sro_n1122;
wire CLOCK_slo__sro_n1123;
wire CLOCK_slo__sro_n1154;
wire CLOCK_slo__sro_n1155;
wire CLOCK_slo__sro_n1156;
wire CLOCK_slo__sro_n1157;
wire CLOCK_slo__sro_n1189;
wire CLOCK_slo__sro_n1190;
wire CLOCK_slo__sro_n1191;
wire CLOCK_slo__sro_n1192;
wire CLOCK_slo__sro_n1193;
wire CLOCK_slo__sro_n1337;
wire CLOCK_slo__sro_n1338;
wire CLOCK_slo__sro_n1339;
wire CLOCK_slo__sro_n1288;
wire CLOCK_slo__sro_n1289;
wire CLOCK_slo__sro_n1290;
wire CLOCK_slo__sro_n1291;


INV_X1 i_36 (.ZN (n_34), .A (p_0[30]));
INV_X1 i_35 (.ZN (n_33), .A (p_1[30]));
INV_X2 i_34 (.ZN (n_32), .A (n_30));
XOR2_X1 i_32 (.Z (p_2[31]), .A (p_0[31]), .B (n_31));
OAI22_X1 i_31 (.ZN (n_0), .A1 (n_34), .A2 (p_1[30]), .B1 (p_0[30]), .B2 (n_33));
XNOR2_X1 i_0 (.ZN (p_2[30]), .A (n_32), .B (n_0));
FA_X1 i_30 (.CO (n_30), .S (p_2[29]), .A (p_0[29]), .B (p_1[29]), .CI (CLOCK_slo__sro_n1190));
INV_X1 CLOCK_slo__sro_c978 (.ZN (CLOCK_slo__sro_n1339), .A (n_30));
FA_X1 i_28 (.CO (n_28), .S (p_2[27]), .A (p_0[27]), .B (p_1[27]), .CI (n_27));
FA_X1 i_27 (.CO (n_27), .S (p_2[26]), .A (p_0[26]), .B (p_1[26]), .CI (n_26));
FA_X1 i_26 (.CO (n_26), .S (p_2[25]), .A (p_0[25]), .B (p_1[25]), .CI (n_25));
FA_X1 i_25 (.CO (n_25), .S (p_2[24]), .A (p_0[24]), .B (p_1[24]), .CI (slo__sro_n155));
NAND2_X1 slo__sro_c168 (.ZN (slo__sro_n243), .A1 (p_1[21]), .A2 (p_0[21]));
FA_X1 i_23 (.CO (n_23), .S (p_2[22]), .A (p_0[22]), .B (p_1[22]), .CI (slo__sro_n241));
INV_X1 slo__sro_c246 (.ZN (slo__sro_n321), .A (n_6));
CLKBUF_X1 slo__L2_c2_c631 (.Z (slo_n883), .A (p_1[13]));
FA_X1 i_20 (.CO (n_20), .S (p_2[19]), .A (p_0[19]), .B (p_1[19]), .CI (slo__sro_n185));
INV_X1 slo__sro_c167 (.ZN (slo__sro_n244), .A (n_21));
FA_X1 i_18 (.CO (n_18), .S (p_2[17]), .A (p_0[17]), .B (p_1[17]), .CI (n_17));
FA_X1 i_17 (.CO (n_17), .S (p_2[16]), .A (p_0[16]), .B (p_1[16]), .CI (n_16));
XNOR2_X2 CLOCK_slo__sro_c772 (.ZN (p_2[4]), .A (CLOCK_slo__sro_n1120), .B (n_4));
NAND2_X1 slo__sro_c543 (.ZN (slo__sro_n756), .A1 (p_1[20]), .A2 (p_0[20]));
INV_X1 CLOCK_slo__sro_c844 (.ZN (CLOCK_slo__sro_n1193), .A (n_28));
FA_X1 i_13 (.CO (n_13), .S (p_2[12]), .A (p_0[12]), .B (p_1[12]), .CI (n_12));
FA_X1 i_11 (.CO (n_11), .S (p_2[10]), .A (p_0[10]), .B (p_1[10]), .CI (n_10));
FA_X1 i_10 (.CO (n_10), .S (p_2[9]), .A (p_0[9]), .B (p_1[9]), .CI (n_9));
FA_X1 i_9 (.CO (n_9), .S (p_2[8]), .A (p_0[8]), .B (p_1[8]), .CI (n_8));
INV_X1 slo__sro_c302 (.ZN (slo__sro_n416), .A (n_14));
INV_X1 slo__sro_c262 (.ZN (slo__sro_n339), .A (slo__n898));
FA_X1 i_6 (.CO (n_6), .S (p_2[5]), .A (p_0[5]), .B (p_1[5]), .CI (n_5));
INV_X2 CLOCK_slo__sro_c804 (.ZN (CLOCK_slo__sro_n1157), .A (n_13));
FA_X1 i_4 (.CO (n_4), .S (p_2[3]), .A (p_0[3]), .B (p_1[3]), .CI (n_3));
FA_X1 i_3 (.CO (n_3), .S (p_2[2]), .A (p_0[2]), .B (p_1[2]), .CI (n_2));
FA_X1 i_2 (.CO (n_2), .S (p_2[1]), .A (p_0[1]), .B (p_1[1]), .CI (n_1));
HA_X1 i_1 (.CO (n_1), .S (p_2[0]), .A (p_0[0]), .B (p_1[0]));
INV_X1 slo__sro_c112 (.ZN (slo__sro_n188), .A (n_18));
NAND2_X1 slo__sro_c113 (.ZN (slo__sro_n187), .A1 (p_1[18]), .A2 (p_0[18]));
NOR2_X1 slo__sro_c114 (.ZN (slo__sro_n186), .A1 (p_1[18]), .A2 (p_0[18]));
OAI21_X1 slo__sro_c115 (.ZN (slo__sro_n185), .A (slo__sro_n187), .B1 (slo__sro_n188), .B2 (slo__sro_n186));
XNOR2_X1 slo__sro_c116 (.ZN (slo__sro_n184), .A (p_1[18]), .B (p_0[18]));
XNOR2_X1 slo__sro_c117 (.ZN (p_2[18]), .A (n_18), .B (slo__sro_n184));
INV_X1 slo__sro_c85 (.ZN (slo__sro_n158), .A (n_23));
NAND2_X1 slo__sro_c86 (.ZN (slo__sro_n157), .A1 (p_1[23]), .A2 (p_0[23]));
NOR2_X1 slo__sro_c87 (.ZN (slo__sro_n156), .A1 (p_1[23]), .A2 (p_0[23]));
OAI21_X1 slo__sro_c88 (.ZN (slo__sro_n155), .A (slo__sro_n157), .B1 (slo__sro_n158), .B2 (slo__sro_n156));
XNOR2_X1 slo__sro_c89 (.ZN (slo__sro_n154), .A (p_1[23]), .B (p_0[23]));
XNOR2_X1 slo__sro_c90 (.ZN (p_2[23]), .A (slo__sro_n154), .B (n_23));
NOR2_X1 slo__sro_c169 (.ZN (slo__sro_n242), .A1 (p_1[21]), .A2 (p_0[21]));
OAI21_X1 slo__sro_c170 (.ZN (slo__sro_n241), .A (slo__sro_n243), .B1 (slo__sro_n242), .B2 (slo__sro_n244));
OAI21_X4 slo__sro_c545 (.ZN (n_21), .A (slo__sro_n756), .B1 (slo__sro_n755), .B2 (slo__sro_n757));
XNOR2_X1 slo__sro_c546 (.ZN (slo__sro_n754), .A (p_1[20]), .B (p_0[20]));
NAND2_X1 slo__sro_c247 (.ZN (slo__sro_n320), .A1 (p_1[6]), .A2 (p_0[6]));
NOR2_X1 slo__sro_c248 (.ZN (slo__sro_n319), .A1 (p_1[6]), .A2 (p_0[6]));
OAI21_X1 slo__sro_c249 (.ZN (slo__sro_n318), .A (slo__sro_n320), .B1 (slo__sro_n321), .B2 (slo__sro_n319));
XNOR2_X1 slo__sro_c250 (.ZN (slo__sro_n317), .A (p_1[6]), .B (p_0[6]));
XNOR2_X1 slo__sro_c251 (.ZN (p_2[6]), .A (n_6), .B (slo__sro_n317));
NAND2_X1 slo__sro_c263 (.ZN (slo__sro_n338), .A1 (p_1[7]), .A2 (p_0[7]));
NOR2_X1 slo__sro_c264 (.ZN (slo__sro_n337), .A1 (p_1[7]), .A2 (p_0[7]));
OAI21_X1 slo__sro_c265 (.ZN (n_8), .A (slo__sro_n338), .B1 (slo__sro_n339), .B2 (slo__sro_n337));
XNOR2_X1 slo__sro_c266 (.ZN (slo__sro_n336), .A (p_1[7]), .B (p_0[7]));
XNOR2_X1 slo__sro_c267 (.ZN (p_2[7]), .A (slo__sro_n336), .B (slo__sro_n318));
NAND2_X1 slo__sro_c303 (.ZN (slo__sro_n415), .A1 (p_1[14]), .A2 (p_0[14]));
NOR2_X1 slo__sro_c304 (.ZN (slo__sro_n414), .A1 (p_1[14]), .A2 (p_0[14]));
OAI21_X1 slo__sro_c305 (.ZN (slo__sro_n413), .A (slo__sro_n415), .B1 (slo__sro_n416), .B2 (slo__sro_n414));
XNOR2_X1 slo__sro_c306 (.ZN (slo__sro_n412), .A (p_1[14]), .B (p_0[14]));
XNOR2_X1 slo__sro_c307 (.ZN (p_2[14]), .A (slo__sro_n412), .B (n_14));
INV_X2 slo__sro_c542 (.ZN (slo__sro_n757), .A (n_20));
NOR2_X1 slo__sro_c544 (.ZN (slo__sro_n755), .A1 (p_1[20]), .A2 (p_0[20]));
XNOR2_X2 slo__mro_c506 (.ZN (slo__mro_n715), .A (n_21), .B (p_0[21]));
XNOR2_X2 slo__mro_c507 (.ZN (p_2[21]), .A (slo__mro_n715), .B (p_1[21]));
XNOR2_X1 slo__sro_c547 (.ZN (p_2[20]), .A (slo__sro_n754), .B (n_20));
OAI21_X1 slo__c638 (.ZN (slo__n898), .A (slo__sro_n320), .B1 (slo__sro_n321), .B2 (slo__sro_n319));
INV_X1 CLOCK_slo__sro_c767 (.ZN (CLOCK_slo__sro_n1123), .A (n_4));
NAND2_X1 CLOCK_slo__sro_c768 (.ZN (CLOCK_slo__sro_n1122), .A1 (p_1[4]), .A2 (p_0[4]));
NOR2_X1 CLOCK_slo__sro_c769 (.ZN (CLOCK_slo__sro_n1121), .A1 (p_1[4]), .A2 (p_0[4]));
OAI21_X1 CLOCK_slo__sro_c770 (.ZN (n_5), .A (CLOCK_slo__sro_n1122), .B1 (CLOCK_slo__sro_n1123), .B2 (CLOCK_slo__sro_n1121));
XNOR2_X2 CLOCK_slo__sro_c771 (.ZN (CLOCK_slo__sro_n1120), .A (p_1[4]), .B (p_0[4]));
INV_X1 slo__sro_c373 (.ZN (slo__sro_n506), .A (slo__sro_n413));
NAND2_X1 slo__sro_c374 (.ZN (slo__sro_n505), .A1 (p_1[15]), .A2 (p_0[15]));
NOR2_X1 slo__sro_c375 (.ZN (slo__sro_n504), .A1 (p_1[15]), .A2 (p_0[15]));
OAI21_X1 slo__sro_c376 (.ZN (n_16), .A (slo__sro_n505), .B1 (slo__sro_n506), .B2 (slo__sro_n504));
XNOR2_X1 slo__sro_c377 (.ZN (slo__sro_n503), .A (p_1[15]), .B (p_0[15]));
XNOR2_X1 slo__sro_c378 (.ZN (p_2[15]), .A (slo__sro_n413), .B (slo__sro_n503));
NAND2_X1 CLOCK_slo__sro_c805 (.ZN (CLOCK_slo__sro_n1156), .A1 (slo_n883), .A2 (p_0[13]));
NOR2_X2 CLOCK_slo__sro_c806 (.ZN (CLOCK_slo__sro_n1155), .A1 (slo_n883), .A2 (p_0[13]));
OAI21_X4 CLOCK_slo__sro_c807 (.ZN (n_14), .A (CLOCK_slo__sro_n1156), .B1 (CLOCK_slo__sro_n1157), .B2 (CLOCK_slo__sro_n1155));
XNOR2_X1 CLOCK_slo__sro_c808 (.ZN (CLOCK_slo__sro_n1154), .A (slo_n883), .B (p_0[13]));
XNOR2_X1 CLOCK_slo__sro_c809 (.ZN (p_2[13]), .A (CLOCK_slo__sro_n1154), .B (n_13));
NAND2_X1 CLOCK_slo__sro_c845 (.ZN (CLOCK_slo__sro_n1192), .A1 (p_1[28]), .A2 (p_0[28]));
NOR2_X1 CLOCK_slo__sro_c846 (.ZN (CLOCK_slo__sro_n1191), .A1 (p_1[28]), .A2 (p_0[28]));
OAI21_X1 CLOCK_slo__sro_c847 (.ZN (CLOCK_slo__sro_n1190), .A (CLOCK_slo__sro_n1192)
    , .B1 (CLOCK_slo__sro_n1193), .B2 (CLOCK_slo__sro_n1191));
XNOR2_X1 CLOCK_slo__sro_c848 (.ZN (CLOCK_slo__sro_n1189), .A (p_1[28]), .B (p_0[28]));
XNOR2_X1 CLOCK_slo__sro_c849 (.ZN (p_2[28]), .A (CLOCK_slo__sro_n1189), .B (n_28));
NOR2_X1 CLOCK_slo__sro_c979 (.ZN (CLOCK_slo__sro_n1338), .A1 (n_33), .A2 (p_0[30]));
NAND2_X1 CLOCK_slo__sro_c980 (.ZN (CLOCK_slo__sro_n1337), .A1 (CLOCK_slo__sro_n1338), .A2 (CLOCK_slo__sro_n1339));
OR2_X1 CLOCK_slo__sro_c981 (.ZN (CLOCK_slo__sro_n1336), .A1 (p_1[30]), .A2 (n_34));
OAI21_X1 CLOCK_slo__sro_c982 (.ZN (n_31), .A (CLOCK_slo__sro_n1337), .B1 (n_32), .B2 (CLOCK_slo__sro_n1336));
INV_X2 CLOCK_slo__sro_c938 (.ZN (CLOCK_slo__sro_n1291), .A (n_11));
NAND2_X1 CLOCK_slo__sro_c939 (.ZN (CLOCK_slo__sro_n1290), .A1 (p_1[11]), .A2 (p_0[11]));
NOR2_X1 CLOCK_slo__sro_c940 (.ZN (CLOCK_slo__sro_n1289), .A1 (p_1[11]), .A2 (p_0[11]));
OAI21_X2 CLOCK_slo__sro_c941 (.ZN (n_12), .A (CLOCK_slo__sro_n1290), .B1 (CLOCK_slo__sro_n1291), .B2 (CLOCK_slo__sro_n1289));
XNOR2_X1 CLOCK_slo__sro_c942 (.ZN (CLOCK_slo__sro_n1288), .A (p_1[11]), .B (p_0[11]));
XNOR2_X1 CLOCK_slo__sro_c943 (.ZN (p_2[11]), .A (n_11), .B (CLOCK_slo__sro_n1288));

endmodule //datapath__0_182

module datapath__0_181 (Multiplier, p_0, p_1);

output [31:0] p_1;
input [31:0] Multiplier;
input [31:0] p_0;
wire slo__n684;
wire slo__sro_n612;
wire n_1;
wire n_2;
wire n_3;
wire n_5;
wire slo__sro_n615;
wire n_7;
wire n_8;
wire n_9;
wire n_10;
wire n_11;
wire n_12;
wire n_13;
wire n_14;
wire n_15;
wire slo__sro_n492;
wire n_17;
wire n_18;
wire slo__sro_n746;
wire n_20;
wire n_21;
wire n_22;
wire n_25;
wire n_26;
wire n_27;
wire n_28;
wire n_30;
wire n_32;
wire n_0;
wire n_34;
wire n_33;
wire spt__n1707;
wire slo__sro_n60;
wire slo__sro_n61;
wire slo__sro_n62;
wire slo__sro_n72;
wire slo__sro_n73;
wire CLOCK_slo__sro_n1121;
wire slo__sro_n75;
wire slo__sro_n85;
wire slo__sro_n86;
wire slo__sro_n87;
wire slo__sro_n88;
wire slo__sro_n98;
wire slo__sro_n99;
wire slo__sro_n100;
wire slo__sro_n101;
wire slo__sro_n113;
wire slo__sro_n114;
wire slo__sro_n115;
wire slo__sro_n116;
wire slo__sro_n117;
wire slo__sro_n144;
wire slo__sro_n145;
wire slo__sro_n146;
wire slo__sro_n147;
wire slo__sro_n148;
wire slo__sro_n164;
wire slo__sro_n165;
wire slo__sro_n178;
wire slo__sro_n179;
wire slo__sro_n180;
wire slo__sro_n181;
wire slo__sro_n182;
wire slo__sro_n493;
wire slo__sro_n494;
wire slo__sro_n613;
wire slo__sro_n614;
wire CLOCK_slo__xsl_n1190;
wire CLOCK_slo__xsl_n1189;
wire slo__sro_n213;
wire slo__sro_n214;
wire slo__sro_n215;
wire slo__sro_n616;
wire slo__sro_n670;
wire slo__sro_n671;
wire slo__sro_n672;
wire slo__sro_n698;
wire slo__sro_n699;
wire slo__sro_n700;
wire slo__sro_n701;
wire slo__mro_n721;
wire slo__sro_n747;
wire slo__sro_n748;
wire slo__sro_n749;
wire slo__sro_n763;
wire slo__sro_n764;
wire slo__sro_n765;
wire slo__sro_n766;
wire slo__sro_n780;
wire slo__sro_n781;
wire slo__sro_n782;
wire slo__sro_n783;
wire slo__sro_n841;
wire CLOCK_slo__sro_n1122;
wire CLOCK_slo__sro_n1123;
wire CLOCK_slo__sro_n1124;
wire CLOCK_slo__sro_n1125;
wire CLOCK_slo__sro_n1142;
wire CLOCK_slo__sro_n1143;
wire CLOCK_slo__sro_n1144;
wire CLOCK_slo__sro_n1145;
wire CLOCK_slo__mro_n1177;
wire CLOCK_slo__mro_n1199;
wire CLOCK_slo__sro_n1285;
wire CLOCK_slo__sro_n1286;
wire CLOCK_slo__sro_n1287;
wire CLOCK_slo__sro_n1288;


INV_X1 i_36 (.ZN (n_34), .A (Multiplier[30]));
INV_X1 i_35 (.ZN (n_33), .A (p_0[30]));
INV_X1 i_34 (.ZN (n_32), .A (n_30));
OAI33_X1 i_33 (.ZN (spt__n1707), .A1 (n_32), .A2 (p_0[30]), .A3 (n_34), .B1 (n_30)
    , .B2 (n_33), .B3 (Multiplier[30]));
XOR2_X1 i_32 (.Z (p_1[31]), .A (Multiplier[31]), .B (spt__n1707));
OAI22_X1 i_31 (.ZN (n_0), .A1 (n_34), .A2 (p_0[30]), .B1 (Multiplier[30]), .B2 (n_33));
XNOR2_X1 i_0 (.ZN (p_1[30]), .A (n_32), .B (n_0));
XNOR2_X1 slo__mro_c529 (.ZN (slo__mro_n721), .A (n_21), .B (Multiplier[21]));
INV_X1 slo__sro_c561 (.ZN (slo__sro_n766), .A (n_17));
INV_X1 slo__sro_c17 (.ZN (slo__sro_n75), .A (n_12));
INV_X1 slo__L1_c494 (.ZN (slo__n684), .A (n_5));
NAND2_X1 slo__sro_c432 (.ZN (slo__sro_n615), .A1 (p_0[23]), .A2 (Multiplier[23]));
FA_X1 i_25 (.CO (n_25), .S (p_1[24]), .A (Multiplier[24]), .B (p_0[24]), .CI (slo__sro_n613));
NAND2_X1 slo__sro_c479 (.ZN (slo__sro_n672), .A1 (p_0[26]), .A2 (Multiplier[26]));
INV_X1 slo__sro_c93 (.ZN (slo__sro_n148), .A (n_18));
INV_X1 slo__sro_c123 (.ZN (slo__sro_n182), .A (n_15));
INV_X1 slo__sro_c64 (.ZN (slo__sro_n117), .A (n_22));
FA_X1 i_20 (.CO (n_20), .S (p_1[19]), .A (Multiplier[19]), .B (p_0[19]), .CI (slo__sro_n145));
INV_X1 slo__sro_c431 (.ZN (slo__sro_n616), .A (slo__sro_n114));
INV_X2 slo__sro_c582 (.ZN (slo__sro_n783), .A (n_11));
FA_X1 i_17 (.CO (n_17), .S (p_1[16]), .A (Multiplier[16]), .B (p_0[16]), .CI (slo__sro_n179));
NAND2_X4 slo__sro_c348 (.ZN (n_26), .A1 (slo__sro_n493), .A2 (slo__sro_n494));
XNOR2_X1 CLOCK_slo__mro_c775 (.ZN (p_1[8]), .A (n_8), .B (slo__sro_n85));
FA_X1 i_14 (.CO (n_14), .S (p_1[13]), .A (Multiplier[13]), .B (p_0[13]), .CI (n_13));
INV_X1 slo__sro_c31 (.ZN (slo__sro_n88), .A (n_8));
INV_X1 CLOCK_slo__sro_c743 (.ZN (CLOCK_slo__sro_n1125), .A (n_3));
FA_X1 i_11 (.CO (n_11), .S (p_1[10]), .A (Multiplier[10]), .B (p_0[10]), .CI (n_10));
INV_X1 slo__sro_c45 (.ZN (slo__sro_n101), .A (n_20));
FA_X1 i_8 (.CO (n_8), .S (p_1[7]), .A (Multiplier[7]), .B (p_0[7]), .CI (n_7));
FA_X1 i_7 (.CO (n_7), .S (p_1[6]), .A (Multiplier[6]), .B (p_0[6]), .CI (slo__sro_n213));
OAI21_X1 slo__sro_c434 (.ZN (slo__sro_n613), .A (slo__sro_n615), .B1 (slo__sro_n616), .B2 (slo__sro_n614));
FA_X1 i_5 (.CO (n_5), .S (p_1[4]), .A (Multiplier[4]), .B (p_0[4]), .CI (CLOCK_slo__sro_n1122));
INV_X1 CLOCK_slo__sro_c761 (.ZN (CLOCK_slo__sro_n1145), .A (n_14));
FA_X1 i_3 (.CO (n_3), .S (p_1[2]), .A (Multiplier[2]), .B (p_0[2]), .CI (n_2));
FA_X1 i_2 (.CO (n_2), .S (p_1[1]), .A (Multiplier[1]), .B (p_0[1]), .CI (n_1));
HA_X1 i_1 (.CO (n_1), .S (p_1[0]), .A (Multiplier[0]), .B (p_0[0]));
INV_X1 slo__sro_c3 (.ZN (slo__sro_n62), .A (n_27));
NAND2_X1 slo__sro_c4 (.ZN (slo__sro_n61), .A1 (p_0[27]), .A2 (Multiplier[27]));
NOR2_X1 slo__sro_c5 (.ZN (slo__sro_n60), .A1 (p_0[27]), .A2 (Multiplier[27]));
OAI21_X1 slo__sro_c6 (.ZN (n_28), .A (slo__sro_n61), .B1 (slo__sro_n60), .B2 (slo__sro_n62));
NOR2_X1 CLOCK_slo__sro_c745 (.ZN (CLOCK_slo__sro_n1123), .A1 (p_0[3]), .A2 (Multiplier[3]));
NOR2_X1 slo__sro_c19 (.ZN (slo__sro_n73), .A1 (p_0[12]), .A2 (Multiplier[12]));
OAI21_X2 slo__sro_c20 (.ZN (n_13), .A (slo__sro_n841), .B1 (slo__sro_n75), .B2 (slo__sro_n73));
XNOR2_X1 slo__sro_c21 (.ZN (slo__sro_n72), .A (p_0[12]), .B (Multiplier[12]));
XNOR2_X1 slo__sro_c22 (.ZN (p_1[12]), .A (slo__sro_n72), .B (n_12));
NAND2_X1 slo__sro_c32 (.ZN (slo__sro_n87), .A1 (p_0[8]), .A2 (Multiplier[8]));
NOR2_X1 slo__sro_c33 (.ZN (slo__sro_n86), .A1 (p_0[8]), .A2 (Multiplier[8]));
OAI21_X2 slo__sro_c34 (.ZN (n_9), .A (slo__sro_n87), .B1 (slo__sro_n88), .B2 (slo__sro_n86));
XNOR2_X1 slo__sro_c35 (.ZN (slo__sro_n85), .A (p_0[8]), .B (Multiplier[8]));
XNOR2_X2 CLOCK_slo__mro_c796 (.ZN (CLOCK_slo__mro_n1177), .A (p_0[5]), .B (Multiplier[5]));
NAND2_X1 slo__sro_c46 (.ZN (slo__sro_n100), .A1 (p_0[20]), .A2 (Multiplier[20]));
NOR2_X1 slo__sro_c47 (.ZN (slo__sro_n99), .A1 (p_0[20]), .A2 (Multiplier[20]));
OAI21_X1 slo__sro_c48 (.ZN (n_21), .A (slo__sro_n100), .B1 (slo__sro_n101), .B2 (slo__sro_n99));
XNOR2_X1 slo__sro_c49 (.ZN (slo__sro_n98), .A (p_0[20]), .B (Multiplier[20]));
XNOR2_X1 slo__sro_c50 (.ZN (p_1[20]), .A (slo__sro_n98), .B (n_20));
NAND2_X1 slo__sro_c65 (.ZN (slo__sro_n116), .A1 (p_0[22]), .A2 (Multiplier[22]));
NOR2_X1 slo__sro_c66 (.ZN (slo__sro_n115), .A1 (p_0[22]), .A2 (Multiplier[22]));
OAI21_X1 slo__sro_c67 (.ZN (slo__sro_n114), .A (slo__sro_n116), .B1 (slo__sro_n117), .B2 (slo__sro_n115));
XNOR2_X2 slo__sro_c68 (.ZN (slo__sro_n113), .A (p_0[22]), .B (Multiplier[22]));
XNOR2_X2 slo__sro_c69 (.ZN (p_1[22]), .A (slo__sro_n113), .B (n_22));
NAND2_X1 slo__sro_c94 (.ZN (slo__sro_n147), .A1 (p_0[18]), .A2 (Multiplier[18]));
NOR2_X1 slo__sro_c95 (.ZN (slo__sro_n146), .A1 (p_0[18]), .A2 (Multiplier[18]));
OAI21_X1 slo__sro_c96 (.ZN (slo__sro_n145), .A (slo__sro_n147), .B1 (slo__sro_n148), .B2 (slo__sro_n146));
XNOR2_X1 slo__sro_c97 (.ZN (slo__sro_n144), .A (p_0[18]), .B (Multiplier[18]));
XNOR2_X1 slo__sro_c98 (.ZN (p_1[18]), .A (slo__sro_n144), .B (n_18));
NAND2_X1 slo__sro_c110 (.ZN (slo__sro_n165), .A1 (p_0[21]), .A2 (Multiplier[21]));
AOI22_X1 slo__sro_c111 (.ZN (slo__sro_n164), .A1 (p_0[21]), .A2 (n_21), .B1 (n_21), .B2 (Multiplier[21]));
NAND2_X1 slo__sro_c112 (.ZN (n_22), .A1 (slo__sro_n165), .A2 (slo__sro_n164));
NAND2_X1 slo__sro_c547 (.ZN (slo__sro_n749), .A1 (n_28), .A2 (Multiplier[28]));
OAI21_X2 slo__sro_c548 (.ZN (slo__sro_n748), .A (p_0[28]), .B1 (n_28), .B2 (Multiplier[28]));
NAND2_X1 slo__sro_c124 (.ZN (slo__sro_n181), .A1 (p_0[15]), .A2 (Multiplier[15]));
NOR2_X1 slo__sro_c125 (.ZN (slo__sro_n180), .A1 (p_0[15]), .A2 (Multiplier[15]));
OAI21_X1 slo__sro_c126 (.ZN (slo__sro_n179), .A (slo__sro_n181), .B1 (slo__sro_n182), .B2 (slo__sro_n180));
XNOR2_X2 slo__sro_c127 (.ZN (slo__sro_n178), .A (p_0[15]), .B (Multiplier[15]));
XNOR2_X2 slo__sro_c128 (.ZN (p_1[15]), .A (slo__sro_n178), .B (n_15));
NAND2_X1 slo__sro_c346 (.ZN (slo__sro_n494), .A1 (p_0[25]), .A2 (Multiplier[25]));
XNOR2_X1 slo__sro_c349 (.ZN (slo__sro_n492), .A (p_0[25]), .B (Multiplier[25]));
XNOR2_X1 slo__sro_c350 (.ZN (p_1[25]), .A (slo__sro_n492), .B (n_25));
NOR2_X1 slo__sro_c433 (.ZN (slo__sro_n614), .A1 (p_0[23]), .A2 (Multiplier[23]));
INV_X1 slo__sro_c509 (.ZN (slo__sro_n701), .A (slo__sro_n747));
NAND2_X1 slo__sro_c153 (.ZN (slo__sro_n215), .A1 (p_0[5]), .A2 (Multiplier[5]));
NOR2_X1 slo__sro_c154 (.ZN (slo__sro_n214), .A1 (p_0[5]), .A2 (Multiplier[5]));
OAI21_X1 slo__sro_c155 (.ZN (slo__sro_n213), .A (slo__sro_n215), .B1 (slo__n684), .B2 (slo__sro_n214));
INV_X1 CLOCK_slo__xsl_c807 (.ZN (CLOCK_slo__xsl_n1190), .A (slo__sro_n114));
INV_X1 CLOCK_slo__xsl_c808 (.ZN (CLOCK_slo__xsl_n1189), .A (CLOCK_slo__xsl_n1190));
XNOR2_X2 slo__sro_c435 (.ZN (slo__sro_n612), .A (p_0[23]), .B (Multiplier[23]));
XNOR2_X2 slo__sro_c436 (.ZN (p_1[23]), .A (slo__sro_n612), .B (CLOCK_slo__xsl_n1189));
AOI22_X2 slo__sro_c480 (.ZN (slo__sro_n671), .A1 (p_0[26]), .A2 (n_26), .B1 (n_26), .B2 (Multiplier[26]));
NAND2_X2 slo__sro_c481 (.ZN (n_27), .A1 (slo__sro_n671), .A2 (slo__sro_n672));
XNOR2_X2 slo__sro_c482 (.ZN (slo__sro_n670), .A (n_26), .B (Multiplier[26]));
XNOR2_X2 slo__sro_c483 (.ZN (p_1[26]), .A (slo__sro_n670), .B (p_0[26]));
NAND2_X1 slo__sro_c510 (.ZN (slo__sro_n700), .A1 (p_0[29]), .A2 (Multiplier[29]));
NOR2_X1 slo__sro_c511 (.ZN (slo__sro_n699), .A1 (p_0[29]), .A2 (Multiplier[29]));
OAI21_X1 slo__sro_c512 (.ZN (n_30), .A (slo__sro_n700), .B1 (slo__sro_n701), .B2 (slo__sro_n699));
XNOR2_X2 slo__sro_c513 (.ZN (slo__sro_n698), .A (p_0[29]), .B (Multiplier[29]));
XNOR2_X1 slo__sro_c514 (.ZN (p_1[29]), .A (slo__sro_n698), .B (slo__sro_n747));
XNOR2_X1 slo__mro_c530 (.ZN (p_1[21]), .A (slo__mro_n721), .B (p_0[21]));
NAND2_X4 slo__sro_c549 (.ZN (slo__sro_n747), .A1 (slo__sro_n748), .A2 (slo__sro_n749));
XNOR2_X2 slo__sro_c550 (.ZN (slo__sro_n746), .A (n_28), .B (Multiplier[28]));
XNOR2_X1 slo__sro_c551 (.ZN (p_1[28]), .A (slo__sro_n746), .B (p_0[28]));
NAND2_X1 slo__sro_c562 (.ZN (slo__sro_n765), .A1 (p_0[17]), .A2 (Multiplier[17]));
NOR2_X1 slo__sro_c563 (.ZN (slo__sro_n764), .A1 (p_0[17]), .A2 (Multiplier[17]));
OAI21_X1 slo__sro_c564 (.ZN (n_18), .A (slo__sro_n765), .B1 (slo__sro_n766), .B2 (slo__sro_n764));
XNOR2_X2 slo__sro_c565 (.ZN (slo__sro_n763), .A (p_0[17]), .B (Multiplier[17]));
XNOR2_X1 slo__sro_c566 (.ZN (p_1[17]), .A (slo__sro_n763), .B (n_17));
NAND2_X1 slo__sro_c583 (.ZN (slo__sro_n782), .A1 (p_0[11]), .A2 (Multiplier[11]));
NOR2_X1 slo__sro_c584 (.ZN (slo__sro_n781), .A1 (p_0[11]), .A2 (Multiplier[11]));
OAI21_X2 slo__sro_c585 (.ZN (n_12), .A (slo__sro_n782), .B1 (slo__sro_n783), .B2 (slo__sro_n781));
XNOR2_X1 slo__sro_c586 (.ZN (slo__sro_n780), .A (p_0[11]), .B (Multiplier[11]));
XNOR2_X1 slo__sro_c587 (.ZN (p_1[11]), .A (slo__sro_n780), .B (n_11));
NAND2_X1 CLOCK_slo__sro_c744 (.ZN (CLOCK_slo__sro_n1124), .A1 (p_0[3]), .A2 (Multiplier[3]));
NAND2_X1 slo__sro_c615 (.ZN (slo__sro_n841), .A1 (p_0[12]), .A2 (Multiplier[12]));
OAI21_X1 CLOCK_slo__sro_c746 (.ZN (CLOCK_slo__sro_n1122), .A (CLOCK_slo__sro_n1124)
    , .B1 (CLOCK_slo__sro_n1123), .B2 (CLOCK_slo__sro_n1125));
XNOR2_X1 CLOCK_slo__sro_c747 (.ZN (CLOCK_slo__sro_n1121), .A (p_0[3]), .B (Multiplier[3]));
XNOR2_X1 CLOCK_slo__sro_c748 (.ZN (p_1[3]), .A (CLOCK_slo__sro_n1121), .B (n_3));
NAND2_X1 CLOCK_slo__sro_c762 (.ZN (CLOCK_slo__sro_n1144), .A1 (p_0[14]), .A2 (Multiplier[14]));
NOR2_X1 CLOCK_slo__sro_c763 (.ZN (CLOCK_slo__sro_n1143), .A1 (p_0[14]), .A2 (Multiplier[14]));
OAI21_X2 CLOCK_slo__sro_c764 (.ZN (n_15), .A (CLOCK_slo__sro_n1144), .B1 (CLOCK_slo__sro_n1145), .B2 (CLOCK_slo__sro_n1143));
XNOR2_X1 CLOCK_slo__sro_c765 (.ZN (CLOCK_slo__sro_n1142), .A (p_0[14]), .B (Multiplier[14]));
XNOR2_X1 CLOCK_slo__sro_c766 (.ZN (p_1[14]), .A (n_14), .B (CLOCK_slo__sro_n1142));
XNOR2_X1 CLOCK_slo__mro_c797 (.ZN (p_1[5]), .A (CLOCK_slo__mro_n1177), .B (n_5));
XNOR2_X2 CLOCK_slo__mro_c815 (.ZN (CLOCK_slo__mro_n1199), .A (n_27), .B (Multiplier[27]));
XNOR2_X2 CLOCK_slo__mro_c816 (.ZN (p_1[27]), .A (CLOCK_slo__mro_n1199), .B (p_0[27]));
INV_X2 CLOCK_slo__sro_c911 (.ZN (CLOCK_slo__sro_n1288), .A (n_9));
NAND2_X1 CLOCK_slo__sro_c912 (.ZN (CLOCK_slo__sro_n1287), .A1 (p_0[9]), .A2 (Multiplier[9]));
NOR2_X1 CLOCK_slo__sro_c913 (.ZN (CLOCK_slo__sro_n1286), .A1 (p_0[9]), .A2 (Multiplier[9]));
OAI21_X1 CLOCK_slo__sro_c914 (.ZN (n_10), .A (CLOCK_slo__sro_n1287), .B1 (CLOCK_slo__sro_n1288), .B2 (CLOCK_slo__sro_n1286));
XNOR2_X1 CLOCK_slo__sro_c915 (.ZN (CLOCK_slo__sro_n1285), .A (p_0[9]), .B (Multiplier[9]));
XNOR2_X1 CLOCK_slo__sro_c916 (.ZN (p_1[9]), .A (CLOCK_slo__sro_n1285), .B (n_9));
OAI21_X2 CLOCK_slo__sro_c944 (.ZN (slo__sro_n493), .A (n_25), .B1 (p_0[25]), .B2 (Multiplier[25]));

endmodule //datapath__0_181

module datapath__0_177 (p_0, p_1, p_2);

output [31:0] p_2;
input [31:0] p_0;
input [31:0] p_1;
wire CLOCK_slo__sro_n1948;
wire slo__sro_n1013;
wire n_1;
wire n_2;
wire n_4;
wire n_5;
wire n_9;
wire n_10;
wire n_11;
wire n_12;
wire slo__sro_n786;
wire n_14;
wire CLOCK_slo__sro_n1947;
wire n_17;
wire n_18;
wire n_19;
wire slo__sro_n215;
wire n_21;
wire CLOCK_slo__sro_n1950;
wire n_23;
wire n_24;
wire n_25;
wire n_26;
wire n_28;
wire n_29;
wire n_30;
wire n_32;
wire n_0;
wire n_34;
wire n_33;
wire n_31;
wire slo__sro_n153;
wire slo__sro_n154;
wire slo__sro_n155;
wire slo__sro_n156;
wire slo__sro_n1010;
wire slo__sro_n212;
wire slo__sro_n213;
wire CLOCK_slo__sro_n1949;
wire slo__sro_n194;
wire slo__sro_n195;
wire slo__sro_n196;
wire slo__sro_n197;
wire slo__sro_n198;
wire slo__sro_n285;
wire slo__sro_n286;
wire slo__sro_n287;
wire slo__sro_n288;
wire slo__sro_n289;
wire slo__mro_n990;
wire slo__sro_n1011;
wire slo__sro_n1012;
wire slo__sro_n784;
wire slo__sro_n785;
wire slo__sro_n429;
wire slo__sro_n430;
wire slo__sro_n431;
wire CLOCK_slo__sro_n1795;
wire slo__sro_n272;
wire slo__sro_n273;
wire slo__sro_n274;
wire slo__sro_n275;
wire slo__sro_n432;
wire slo__sro_n433;
wire slo__sro_n620;
wire slo__sro_n621;
wire slo__sro_n622;
wire slo__sro_n623;
wire slo__sro_n787;
wire slo__sro_n1014;
wire CLOCK_slo__sro_n1530;
wire CLOCK_slo__sro_n1531;
wire CLOCK_slo__sro_n1532;
wire CLOCK_slo__sro_n1533;
wire CLOCK_slo__sro_n1534;
wire slo__sro_n1073;
wire slo__sro_n1074;
wire slo__sro_n1075;
wire slo__sro_n1076;
wire slo__sro_n1077;
wire CLOCK_slo__sro_n1602;
wire CLOCK_slo__sro_n1603;
wire CLOCK_slo__sro_n1604;
wire CLOCK_slo__sro_n1605;
wire CLOCK_slo__sro_n1606;
wire CLOCK_slo__sro_n1653;
wire CLOCK_slo__sro_n1654;
wire CLOCK_slo__sro_n1655;
wire CLOCK_slo__sro_n1656;
wire CLOCK_slo__sro_n1666;
wire CLOCK_slo__sro_n1667;
wire CLOCK_slo__sro_n1668;
wire CLOCK_slo__sro_n1669;


INV_X1 i_36 (.ZN (n_34), .A (p_0[30]));
INV_X1 i_35 (.ZN (n_33), .A (p_1[30]));
INV_X1 i_34 (.ZN (n_32), .A (n_30));
OAI33_X1 i_33 (.ZN (n_31), .A1 (n_32), .A2 (p_1[30]), .A3 (n_34), .B1 (n_30), .B2 (n_33), .B3 (p_0[30]));
XOR2_X1 i_32 (.Z (p_2[31]), .A (p_0[31]), .B (n_31));
OAI22_X1 i_31 (.ZN (n_0), .A1 (n_34), .A2 (p_1[30]), .B1 (p_0[30]), .B2 (n_33));
XNOR2_X1 i_0 (.ZN (p_2[30]), .A (n_32), .B (n_0));
XNOR2_X1 slo__sro_c722 (.ZN (p_2[26]), .A (slo__sro_n1010), .B (n_26));
FA_X1 i_29 (.CO (n_29), .S (p_2[28]), .A (p_0[28]), .B (p_1[28]), .CI (n_28));
FA_X1 i_28 (.CO (n_28), .S (p_2[27]), .A (p_0[27]), .B (p_1[27]), .CI (slo__sro_n1011));
INV_X1 CLOCK_slo__sro_c982 (.ZN (CLOCK_slo__sro_n1534), .A (n_2));
FA_X1 i_26 (.CO (n_26), .S (p_2[25]), .A (p_0[25]), .B (p_1[25]), .CI (n_25));
FA_X1 i_25 (.CO (n_25), .S (p_2[24]), .A (p_0[24]), .B (p_1[24]), .CI (n_24));
INV_X1 slo__sro_c141 (.ZN (slo__sro_n215), .A (n_5));
FA_X1 i_23 (.CO (n_23), .S (p_2[22]), .A (p_0[22]), .B (p_1[22]), .CI (CLOCK_slo__sro_n1667));
XNOR2_X2 CLOCK_slo__sro_c1376 (.ZN (p_2[6]), .A (CLOCK_slo__sro_n1947), .B (slo__sro_n212));
NAND2_X1 CLOCK_slo__sro_c1120 (.ZN (CLOCK_slo__sro_n1669), .A1 (n_21), .A2 (p_0[21]));
NAND2_X1 slo__sro_c211 (.ZN (slo__sro_n288), .A1 (p_1[7]), .A2 (p_0[7]));
FA_X1 i_19 (.CO (n_19), .S (p_2[18]), .A (p_0[18]), .B (p_1[18]), .CI (n_18));
XNOR2_X1 slo__sro_c603 (.ZN (p_2[29]), .A (n_29), .B (slo__sro_n784));
FA_X1 i_17 (.CO (n_17), .S (p_2[16]), .A (p_0[16]), .B (p_1[16]), .CI (slo__sro_n1074));
NAND2_X1 CLOCK_slo__sro_c1372 (.ZN (CLOCK_slo__sro_n1950), .A1 (p_1[6]), .A2 (p_0[6]));
NAND2_X1 CLOCK_slo__sro_c1106 (.ZN (CLOCK_slo__sro_n1656), .A1 (p_1[20]), .A2 (p_0[20]));
XNOR2_X1 slo__sro_c305 (.ZN (slo__sro_n429), .A (p_1[12]), .B (p_0[12]));
OAI21_X1 slo__sro_c601 (.ZN (n_30), .A (slo__sro_n786), .B1 (slo__sro_n787), .B2 (slo__sro_n785));
FA_X1 i_12 (.CO (n_12), .S (p_2[11]), .A (p_0[11]), .B (p_1[11]), .CI (n_11));
FA_X1 i_11 (.CO (n_11), .S (p_2[10]), .A (p_0[10]), .B (p_1[10]), .CI (n_10));
FA_X1 i_10 (.CO (n_10), .S (p_2[9]), .A (p_0[9]), .B (p_1[9]), .CI (n_9));
FA_X1 i_9 (.CO (n_9), .S (p_2[8]), .A (p_0[8]), .B (p_1[8]), .CI (slo__sro_n286));
NAND2_X1 CLOCK_slo__sro_c1374 (.ZN (CLOCK_slo__sro_n1948), .A1 (CLOCK_slo__sro_n1949), .A2 (CLOCK_slo__sro_n1950));
INV_X1 slo__sro_c210 (.ZN (slo__sro_n289), .A (CLOCK_slo__sro_n1948));
FA_X1 i_5 (.CO (n_5), .S (p_2[4]), .A (p_0[4]), .B (p_1[4]), .CI (n_4));
FA_X1 i_4 (.CO (n_4), .S (p_2[3]), .A (p_0[3]), .B (p_1[3]), .CI (CLOCK_slo__sro_n1531));
OAI21_X1 CLOCK_slo__sro_c1373 (.ZN (CLOCK_slo__sro_n1949), .A (slo__sro_n212), .B1 (p_1[6]), .B2 (p_0[6]));
FA_X1 i_2 (.CO (n_2), .S (p_2[1]), .A (p_0[1]), .B (p_1[1]), .CI (n_1));
HA_X1 i_1 (.CO (n_1), .S (p_2[0]), .A (p_0[0]), .B (p_1[0]));
INV_X1 slo__sro_c85 (.ZN (slo__sro_n156), .A (n_23));
NAND2_X1 slo__sro_c86 (.ZN (slo__sro_n155), .A1 (p_1[23]), .A2 (p_0[23]));
NOR2_X1 slo__sro_c87 (.ZN (slo__sro_n154), .A1 (p_1[23]), .A2 (p_0[23]));
OAI21_X1 slo__sro_c88 (.ZN (n_24), .A (slo__sro_n155), .B1 (slo__sro_n156), .B2 (slo__sro_n154));
XNOR2_X2 slo__sro_c89 (.ZN (slo__sro_n153), .A (p_1[23]), .B (p_0[23]));
XNOR2_X1 slo__sro_c90 (.ZN (p_2[23]), .A (slo__sro_n153), .B (n_23));
NOR2_X1 slo__sro_c143 (.ZN (slo__sro_n213), .A1 (p_1[5]), .A2 (p_0[5]));
XNOR2_X1 CLOCK_slo__sro_c1168 (.ZN (p_2[13]), .A (slo__sro_n430), .B (slo__sro_n272));
INV_X1 slo__sro_c717 (.ZN (slo__sro_n1014), .A (n_26));
NAND2_X1 slo__sro_c718 (.ZN (slo__sro_n1013), .A1 (p_1[26]), .A2 (p_0[26]));
INV_X1 slo__sro_c127 (.ZN (slo__sro_n198), .A (n_19));
NAND2_X1 slo__sro_c128 (.ZN (slo__sro_n197), .A1 (p_1[19]), .A2 (p_0[19]));
NOR2_X1 slo__sro_c129 (.ZN (slo__sro_n196), .A1 (p_1[19]), .A2 (p_0[19]));
OAI21_X1 slo__sro_c130 (.ZN (slo__sro_n195), .A (slo__sro_n197), .B1 (slo__sro_n198), .B2 (slo__sro_n196));
XNOR2_X1 slo__sro_c131 (.ZN (slo__sro_n194), .A (p_1[19]), .B (p_0[19]));
XNOR2_X1 slo__sro_c132 (.ZN (p_2[19]), .A (slo__sro_n194), .B (n_19));
NOR2_X1 slo__sro_c212 (.ZN (slo__sro_n287), .A1 (p_1[7]), .A2 (p_0[7]));
OAI21_X1 slo__sro_c213 (.ZN (slo__sro_n286), .A (slo__sro_n288), .B1 (slo__sro_n289), .B2 (slo__sro_n287));
XNOR2_X1 slo__sro_c214 (.ZN (slo__sro_n285), .A (p_1[7]), .B (p_0[7]));
XNOR2_X1 slo__sro_c215 (.ZN (p_2[7]), .A (slo__sro_n285), .B (CLOCK_slo__sro_n1948));
XNOR2_X2 slo__mro_c707 (.ZN (slo__mro_n990), .A (n_5), .B (p_0[5]));
XNOR2_X1 slo__mro_c708 (.ZN (p_2[5]), .A (slo__mro_n990), .B (p_1[5]));
NOR2_X1 slo__sro_c719 (.ZN (slo__sro_n1012), .A1 (p_1[26]), .A2 (p_0[26]));
OAI21_X1 slo__sro_c720 (.ZN (slo__sro_n1011), .A (slo__sro_n1013), .B1 (slo__sro_n1012), .B2 (slo__sro_n1014));
XNOR2_X1 slo__sro_c721 (.ZN (slo__sro_n1010), .A (p_1[26]), .B (p_0[26]));
INV_X1 slo__sro_c598 (.ZN (slo__sro_n787), .A (n_29));
NAND2_X1 slo__sro_c599 (.ZN (slo__sro_n786), .A1 (p_1[29]), .A2 (p_0[29]));
NOR2_X1 slo__sro_c600 (.ZN (slo__sro_n785), .A1 (p_1[29]), .A2 (p_0[29]));
INV_X1 slo__sro_c301 (.ZN (slo__sro_n433), .A (n_12));
NAND2_X1 slo__sro_c302 (.ZN (slo__sro_n432), .A1 (p_1[12]), .A2 (p_0[12]));
NOR2_X1 slo__sro_c303 (.ZN (slo__sro_n431), .A1 (p_1[12]), .A2 (p_0[12]));
OAI21_X1 slo__sro_c304 (.ZN (slo__sro_n430), .A (slo__sro_n432), .B1 (slo__sro_n433), .B2 (slo__sro_n431));
INV_X1 slo__sro_c196 (.ZN (slo__sro_n275), .A (slo__sro_n430));
NAND2_X1 slo__sro_c197 (.ZN (slo__sro_n274), .A1 (p_1[13]), .A2 (p_0[13]));
NOR2_X1 slo__sro_c198 (.ZN (slo__sro_n273), .A1 (p_1[13]), .A2 (p_0[13]));
OAI21_X2 slo__sro_c199 (.ZN (n_14), .A (slo__sro_n274), .B1 (slo__sro_n275), .B2 (slo__sro_n273));
XNOR2_X1 slo__sro_c200 (.ZN (slo__sro_n272), .A (p_1[13]), .B (p_0[13]));
XNOR2_X2 CLOCK_slo__sro_c1375 (.ZN (CLOCK_slo__sro_n1947), .A (p_1[6]), .B (p_0[6]));
XNOR2_X1 slo__sro_c306 (.ZN (p_2[12]), .A (slo__sro_n429), .B (n_12));
XNOR2_X1 slo__sro_c602 (.ZN (slo__sro_n784), .A (p_1[29]), .B (p_0[29]));
INV_X1 slo__sro_c457 (.ZN (slo__sro_n623), .A (n_17));
NAND2_X1 slo__sro_c458 (.ZN (slo__sro_n622), .A1 (p_1[17]), .A2 (p_0[17]));
NOR2_X1 slo__sro_c459 (.ZN (slo__sro_n621), .A1 (p_1[17]), .A2 (p_0[17]));
OAI21_X1 slo__sro_c460 (.ZN (n_18), .A (slo__sro_n622), .B1 (slo__sro_n623), .B2 (slo__sro_n621));
XNOR2_X1 slo__sro_c461 (.ZN (slo__sro_n620), .A (p_1[17]), .B (p_0[17]));
XNOR2_X1 slo__sro_c462 (.ZN (p_2[17]), .A (slo__sro_n620), .B (n_17));
NAND2_X1 CLOCK_slo__sro_c983 (.ZN (CLOCK_slo__sro_n1533), .A1 (p_1[2]), .A2 (p_0[2]));
NOR2_X1 CLOCK_slo__sro_c984 (.ZN (CLOCK_slo__sro_n1532), .A1 (p_1[2]), .A2 (p_0[2]));
OAI21_X1 CLOCK_slo__sro_c985 (.ZN (CLOCK_slo__sro_n1531), .A (CLOCK_slo__sro_n1533)
    , .B1 (CLOCK_slo__sro_n1532), .B2 (CLOCK_slo__sro_n1534));
XNOR2_X2 CLOCK_slo__sro_c986 (.ZN (CLOCK_slo__sro_n1530), .A (p_1[2]), .B (p_0[2]));
XNOR2_X1 CLOCK_slo__sro_c987 (.ZN (p_2[2]), .A (CLOCK_slo__sro_n1530), .B (n_2));
INV_X1 slo__sro_c774 (.ZN (slo__sro_n1077), .A (CLOCK_slo__sro_n1603));
NAND2_X1 slo__sro_c775 (.ZN (slo__sro_n1076), .A1 (p_1[15]), .A2 (p_0[15]));
NOR2_X1 slo__sro_c776 (.ZN (slo__sro_n1075), .A1 (p_1[15]), .A2 (p_0[15]));
OAI21_X1 slo__sro_c777 (.ZN (slo__sro_n1074), .A (slo__sro_n1076), .B1 (slo__sro_n1077), .B2 (slo__sro_n1075));
XNOR2_X1 slo__sro_c778 (.ZN (slo__sro_n1073), .A (p_1[15]), .B (p_0[15]));
XNOR2_X1 slo__sro_c779 (.ZN (p_2[15]), .A (slo__sro_n1073), .B (CLOCK_slo__sro_n1603));
INV_X1 CLOCK_slo__sro_c1062 (.ZN (CLOCK_slo__sro_n1606), .A (n_14));
NAND2_X1 CLOCK_slo__sro_c1063 (.ZN (CLOCK_slo__sro_n1605), .A1 (p_1[14]), .A2 (p_0[14]));
NOR2_X1 CLOCK_slo__sro_c1064 (.ZN (CLOCK_slo__sro_n1604), .A1 (p_1[14]), .A2 (p_0[14]));
OAI21_X2 CLOCK_slo__sro_c1065 (.ZN (CLOCK_slo__sro_n1603), .A (CLOCK_slo__sro_n1605)
    , .B1 (CLOCK_slo__sro_n1606), .B2 (CLOCK_slo__sro_n1604));
XNOR2_X1 CLOCK_slo__sro_c1066 (.ZN (CLOCK_slo__sro_n1602), .A (p_1[14]), .B (p_0[14]));
XNOR2_X1 CLOCK_slo__sro_c1067 (.ZN (p_2[14]), .A (CLOCK_slo__sro_n1602), .B (n_14));
NAND2_X1 CLOCK_slo__sro_c1107 (.ZN (CLOCK_slo__sro_n1655), .A1 (slo__sro_n195), .A2 (p_0[20]));
NAND2_X1 CLOCK_slo__sro_c1108 (.ZN (CLOCK_slo__sro_n1654), .A1 (slo__sro_n195), .A2 (p_1[20]));
NAND3_X1 CLOCK_slo__sro_c1109 (.ZN (n_21), .A1 (CLOCK_slo__sro_n1655), .A2 (CLOCK_slo__sro_n1654), .A3 (CLOCK_slo__sro_n1656));
XNOR2_X1 CLOCK_slo__sro_c1110 (.ZN (CLOCK_slo__sro_n1653), .A (p_1[20]), .B (p_0[20]));
XNOR2_X1 CLOCK_slo__sro_c1111 (.ZN (p_2[20]), .A (CLOCK_slo__sro_n1653), .B (slo__sro_n195));
OAI21_X1 CLOCK_slo__sro_c1121 (.ZN (CLOCK_slo__sro_n1668), .A (p_1[21]), .B1 (n_21), .B2 (p_0[21]));
NAND2_X1 CLOCK_slo__sro_c1122 (.ZN (CLOCK_slo__sro_n1667), .A1 (CLOCK_slo__sro_n1668), .A2 (CLOCK_slo__sro_n1669));
XNOR2_X1 CLOCK_slo__sro_c1123 (.ZN (CLOCK_slo__sro_n1666), .A (n_21), .B (p_0[21]));
XNOR2_X1 CLOCK_slo__sro_c1124 (.ZN (p_2[21]), .A (CLOCK_slo__sro_n1666), .B (p_1[21]));
OAI21_X1 CLOCK_slo__sro_c1158 (.ZN (slo__sro_n212), .A (CLOCK_slo__sro_n1795), .B1 (slo__sro_n213), .B2 (slo__sro_n215));
NAND2_X1 CLOCK_slo__sro_c1220 (.ZN (CLOCK_slo__sro_n1795), .A1 (p_1[5]), .A2 (p_0[5]));

endmodule //datapath__0_177

module datapath__0_176 (Multiplier, p_0, p_1);

output [31:0] p_1;
input [31:0] Multiplier;
input [31:0] p_0;
wire CLOCK_slo__sro_n1618;
wire slo__mro_n1013;
wire n_1;
wire n_2;
wire n_3;
wire n_4;
wire n_5;
wire n_7;
wire n_9;
wire n_11;
wire n_12;
wire n_13;
wire n_14;
wire n_15;
wire n_16;
wire n_17;
wire n_18;
wire n_19;
wire n_20;
wire n_21;
wire n_22;
wire n_24;
wire n_25;
wire n_28;
wire n_30;
wire n_32;
wire n_0;
wire n_34;
wire n_33;
wire n_31;
wire slo__sro_n61;
wire slo__sro_n62;
wire slo__sro_n63;
wire slo__sro_n64;
wire slo__sro_n74;
wire slo__sro_n75;
wire slo__sro_n76;
wire slo__sro_n77;
wire slo__sro_n153;
wire slo__sro_n154;
wire slo__sro_n155;
wire slo__sro_n156;
wire CLOCK_slo__sro_n1597;
wire slo__sro_n184;
wire slo__sro_n185;
wire slo__sro_n186;
wire slo__sro_n198;
wire slo__sro_n199;
wire slo__sro_n200;
wire slo__sro_n201;
wire slo__sro_n228;
wire slo__sro_n229;
wire slo__sro_n230;
wire slo__sro_n231;
wire slo__sro_n232;
wire slo__sro_n245;
wire slo__sro_n247;
wire slo__sro_n254;
wire slo__sro_n260;
wire slo__sro_n261;
wire slo__sro_n262;
wire slo__sro_n263;
wire CLOCK_slo__sro_n1683;
wire slo__sro_n280;
wire slo__sro_n281;
wire slo__sro_n282;
wire slo__sro_n309;
wire slo__sro_n310;
wire slo__sro_n311;
wire slo__sro_n312;
wire slo__sro_n324;
wire slo__sro_n325;
wire slo__sro_n326;
wire slo__sro_n327;
wire slo__sro_n328;
wire slo__sro_n496;
wire slo__sro_n497;
wire slo__sro_n498;
wire slo__sro_n499;
wire slo__sro_n753;
wire slo__sro_n537;
wire slo__sro_n538;
wire slo__sro_n539;
wire slo__sro_n754;
wire CLOCK_slo__sro_n1568;
wire slo__sro_n755;
wire slo__sro_n756;
wire CLOCK_slo__sro_n1565;
wire CLOCK_slo__sro_n1566;
wire CLOCK_slo__sro_n1567;
wire CLOCK_slo__sro_n1569;
wire CLOCK_slo__mro_n1584;
wire CLOCK_slo__sro_n1598;
wire CLOCK_slo__sro_n1599;
wire CLOCK_slo__sro_n1600;
wire CLOCK_slo__sro_n1619;
wire CLOCK_slo__sro_n1620;
wire CLOCK_slo__sro_n1621;
wire CLOCK_slo__sro_n1622;
wire CLOCK_slo__sro_n1623;
wire CLOCK_slo__xsl_n1652;
wire CLOCK_slo__sro_n1682;
wire CLOCK_slo__sro_n1684;
wire CLOCK_slo__sro_n1685;
wire CLOCK_slo__mro_n1721;
wire CLOCK_slo__mro_n1722;
wire CLOCK_slo__mro_n1723;
wire CLOCK_slo__sro_n1860;


INV_X1 i_36 (.ZN (n_34), .A (Multiplier[30]));
INV_X1 i_35 (.ZN (n_33), .A (p_0[30]));
INV_X1 i_34 (.ZN (n_32), .A (n_30));
NAND2_X1 CLOCK_slo__sro_c1102 (.ZN (CLOCK_slo__sro_n1685), .A1 (CLOCK_slo__sro_n1860), .A2 (Multiplier[26]));
XOR2_X1 i_32 (.Z (p_1[31]), .A (Multiplier[31]), .B (n_31));
OAI22_X1 i_31 (.ZN (n_0), .A1 (n_34), .A2 (p_0[30]), .B1 (Multiplier[30]), .B2 (n_33));
XNOR2_X1 i_0 (.ZN (p_1[30]), .A (n_32), .B (n_0));
FA_X1 i_30 (.CO (n_30), .S (p_1[29]), .A (Multiplier[29]), .B (p_0[29]), .CI (CLOCK_slo__sro_n1566));
XNOR2_X2 CLOCK_slo__mro_c991 (.ZN (CLOCK_slo__mro_n1584), .A (n_22), .B (Multiplier[22]));
INV_X1 CLOCK_slo__sro_c1021 (.ZN (CLOCK_slo__sro_n1623), .A (n_34));
INV_X1 CLOCK_slo__mro_c1141 (.ZN (slo__mro_n1013), .A (Multiplier[8]));
INV_X2 slo__sro_c166 (.ZN (slo__sro_n232), .A (n_7));
FA_X1 i_25 (.CO (n_25), .S (p_1[24]), .A (Multiplier[24]), .B (p_0[24]), .CI (n_24));
INV_X1 slo__sro_c98 (.ZN (slo__sro_n156), .A (n_19));
INV_X1 slo__sro_c139 (.ZN (slo__sro_n201), .A (n_25));
INV_X1 slo__sro_c548 (.ZN (slo__sro_n756), .A (n_16));
OAI21_X1 slo__sro_c192 (.ZN (slo__sro_n254), .A (n_20), .B1 (p_0[20]), .B2 (Multiplier[20]));
NAND2_X1 slo__sro_c127 (.ZN (slo__sro_n186), .A1 (p_0[22]), .A2 (Multiplier[22]));
FA_X1 i_19 (.CO (n_19), .S (p_1[18]), .A (Multiplier[18]), .B (p_0[18]), .CI (n_18));
INV_X1 slo__sro_c253 (.ZN (slo__sro_n328), .A (p_0[5]));
FA_X1 i_16 (.CO (n_16), .S (p_1[15]), .A (Multiplier[15]), .B (p_0[15]), .CI (n_15));
INV_X1 slo__sro_c17 (.ZN (slo__sro_n77), .A (slo__sro_n184));
FA_X1 i_14 (.CO (n_14), .S (p_1[13]), .A (Multiplier[13]), .B (p_0[13]), .CI (n_13));
NOR2_X1 slo__sro_c550 (.ZN (slo__sro_n754), .A1 (p_0[16]), .A2 (Multiplier[16]));
FA_X1 i_12 (.CO (n_12), .S (p_1[11]), .A (Multiplier[11]), .B (p_0[11]), .CI (n_11));
FA_X1 i_11 (.CO (n_11), .S (p_1[10]), .A (Multiplier[10]), .B (p_0[10]), .CI (slo__sro_n261));
NAND2_X1 slo__sro_c212 (.ZN (slo__sro_n282), .A1 (p_0[8]), .A2 (Multiplier[8]));
INV_X2 slo__sro_c239 (.ZN (slo__sro_n312), .A (n_17));
NAND2_X1 slo__sro_c180 (.ZN (slo__sro_n247), .A1 (p_0[20]), .A2 (Multiplier[20]));
FA_X1 i_7 (.CO (n_7), .S (p_1[6]), .A (Multiplier[6]), .B (p_0[6]), .CI (slo__sro_n325));
INV_X1 slo__sro_c351 (.ZN (slo__sro_n499), .A (n_12));
FA_X1 i_5 (.CO (n_5), .S (p_1[4]), .A (Multiplier[4]), .B (p_0[4]), .CI (n_4));
FA_X1 i_4 (.CO (n_4), .S (p_1[3]), .A (Multiplier[3]), .B (p_0[3]), .CI (n_3));
FA_X1 i_3 (.CO (n_3), .S (p_1[2]), .A (Multiplier[2]), .B (p_0[2]), .CI (n_2));
FA_X1 i_2 (.CO (n_2), .S (p_1[1]), .A (Multiplier[1]), .B (p_0[1]), .CI (n_1));
HA_X1 i_1 (.CO (n_1), .S (p_1[0]), .A (Multiplier[0]), .B (p_0[0]));
INV_X1 slo__sro_c3 (.ZN (slo__sro_n64), .A (n_14));
NAND2_X1 slo__sro_c4 (.ZN (slo__sro_n63), .A1 (p_0[14]), .A2 (Multiplier[14]));
NOR2_X1 slo__sro_c5 (.ZN (slo__sro_n62), .A1 (p_0[14]), .A2 (Multiplier[14]));
OAI21_X1 slo__sro_c6 (.ZN (n_15), .A (slo__sro_n63), .B1 (slo__sro_n64), .B2 (slo__sro_n62));
XNOR2_X1 slo__sro_c7 (.ZN (slo__sro_n61), .A (p_0[14]), .B (Multiplier[14]));
XNOR2_X1 slo__sro_c8 (.ZN (p_1[14]), .A (n_14), .B (slo__sro_n61));
NAND2_X1 slo__sro_c18 (.ZN (slo__sro_n76), .A1 (p_0[23]), .A2 (Multiplier[23]));
NOR2_X2 slo__sro_c19 (.ZN (slo__sro_n75), .A1 (p_0[23]), .A2 (Multiplier[23]));
XNOR2_X1 slo__sro_c21 (.ZN (slo__sro_n74), .A (p_0[23]), .B (Multiplier[23]));
XNOR2_X2 slo__sro_c22 (.ZN (p_1[23]), .A (slo__sro_n74), .B (slo__sro_n184));
NAND2_X1 slo__sro_c99 (.ZN (slo__sro_n155), .A1 (p_0[19]), .A2 (Multiplier[19]));
NOR2_X1 slo__sro_c100 (.ZN (slo__sro_n154), .A1 (p_0[19]), .A2 (Multiplier[19]));
OAI21_X2 slo__sro_c101 (.ZN (n_20), .A (slo__sro_n155), .B1 (slo__sro_n156), .B2 (slo__sro_n154));
XNOR2_X1 slo__sro_c102 (.ZN (slo__sro_n153), .A (p_0[19]), .B (Multiplier[19]));
XNOR2_X1 slo__sro_c103 (.ZN (p_1[19]), .A (slo__sro_n153), .B (n_19));
OAI21_X1 slo__sro_c128 (.ZN (slo__sro_n185), .A (n_22), .B1 (p_0[22]), .B2 (Multiplier[22]));
NAND2_X1 slo__sro_c129 (.ZN (slo__sro_n184), .A1 (slo__sro_n185), .A2 (slo__sro_n186));
INV_X1 CLOCK_slo__sro_c1001 (.ZN (CLOCK_slo__sro_n1600), .A (CLOCK_slo__sro_n1683));
NAND2_X1 CLOCK_slo__sro_c1002 (.ZN (CLOCK_slo__sro_n1599), .A1 (p_0[27]), .A2 (Multiplier[27]));
NAND2_X1 slo__sro_c140 (.ZN (slo__sro_n200), .A1 (p_0[25]), .A2 (Multiplier[25]));
NOR2_X1 slo__sro_c141 (.ZN (slo__sro_n199), .A1 (p_0[25]), .A2 (Multiplier[25]));
XNOR2_X2 slo__sro_c143 (.ZN (slo__sro_n198), .A (p_0[25]), .B (Multiplier[25]));
XNOR2_X2 slo__sro_c144 (.ZN (p_1[25]), .A (slo__sro_n198), .B (n_25));
NAND2_X1 slo__sro_c167 (.ZN (slo__sro_n231), .A1 (p_0[7]), .A2 (Multiplier[7]));
NOR2_X1 slo__sro_c168 (.ZN (slo__sro_n230), .A1 (p_0[7]), .A2 (Multiplier[7]));
OAI21_X2 slo__sro_c169 (.ZN (slo__sro_n229), .A (slo__sro_n231), .B1 (slo__sro_n232), .B2 (slo__sro_n230));
XNOR2_X1 slo__sro_c170 (.ZN (slo__sro_n228), .A (p_0[7]), .B (Multiplier[7]));
XNOR2_X1 slo__sro_c171 (.ZN (p_1[7]), .A (slo__sro_n228), .B (n_7));
XNOR2_X1 CLOCK_slo__sro_c1106 (.ZN (p_1[26]), .A (CLOCK_slo__sro_n1682), .B (p_0[26]));
NAND2_X1 slo__sro_c182 (.ZN (n_21), .A1 (slo__sro_n247), .A2 (slo__sro_n254));
XNOR2_X1 slo__sro_c183 (.ZN (slo__sro_n245), .A (n_20), .B (Multiplier[20]));
NAND2_X1 slo__sro_c197 (.ZN (slo__sro_n263), .A1 (p_0[9]), .A2 (Multiplier[9]));
NOR2_X1 slo__sro_c198 (.ZN (slo__sro_n262), .A1 (p_0[9]), .A2 (Multiplier[9]));
OAI21_X1 slo__sro_c199 (.ZN (slo__sro_n261), .A (slo__sro_n263), .B1 (slo__sro_n262), .B2 (n_9));
XNOR2_X1 slo__sro_c200 (.ZN (slo__sro_n260), .A (p_0[9]), .B (Multiplier[9]));
XNOR2_X1 slo__sro_c201 (.ZN (p_1[9]), .A (slo__sro_n260), .B (CLOCK_slo__xsl_n1652));
NAND2_X2 slo__sro_c213 (.ZN (slo__sro_n281), .A1 (slo__sro_n229), .A2 (Multiplier[8]));
NAND2_X1 slo__sro_c214 (.ZN (slo__sro_n280), .A1 (p_0[8]), .A2 (slo__sro_n229));
OAI21_X1 CLOCK_slo__mro_c1142 (.ZN (CLOCK_slo__mro_n1723), .A (slo__sro_n231), .B1 (slo__sro_n232), .B2 (slo__sro_n230));
INV_X1 CLOCK_slo__sro_c975 (.ZN (CLOCK_slo__sro_n1569), .A (n_28));
NAND2_X1 slo__sro_c240 (.ZN (slo__sro_n311), .A1 (p_0[17]), .A2 (Multiplier[17]));
NOR2_X1 slo__sro_c241 (.ZN (slo__sro_n310), .A1 (p_0[17]), .A2 (Multiplier[17]));
OAI21_X1 slo__sro_c242 (.ZN (n_18), .A (slo__sro_n311), .B1 (slo__sro_n312), .B2 (slo__sro_n310));
XNOR2_X1 slo__sro_c243 (.ZN (slo__sro_n309), .A (p_0[17]), .B (Multiplier[17]));
XNOR2_X1 slo__sro_c244 (.ZN (p_1[17]), .A (slo__sro_n309), .B (n_17));
NAND2_X1 slo__sro_c254 (.ZN (slo__sro_n327), .A1 (n_5), .A2 (Multiplier[5]));
NOR2_X1 slo__sro_c255 (.ZN (slo__sro_n326), .A1 (n_5), .A2 (Multiplier[5]));
OAI21_X1 slo__sro_c256 (.ZN (slo__sro_n325), .A (slo__sro_n327), .B1 (slo__sro_n326), .B2 (slo__sro_n328));
XNOR2_X2 slo__sro_c257 (.ZN (slo__sro_n324), .A (n_5), .B (Multiplier[5]));
XNOR2_X1 slo__sro_c258 (.ZN (p_1[5]), .A (slo__sro_n324), .B (p_0[5]));
NAND2_X1 slo__sro_c352 (.ZN (slo__sro_n498), .A1 (p_0[12]), .A2 (Multiplier[12]));
NOR2_X1 slo__sro_c353 (.ZN (slo__sro_n497), .A1 (p_0[12]), .A2 (Multiplier[12]));
OAI21_X1 slo__sro_c354 (.ZN (n_13), .A (slo__sro_n498), .B1 (slo__sro_n499), .B2 (slo__sro_n497));
XNOR2_X1 slo__sro_c355 (.ZN (slo__sro_n496), .A (p_0[12]), .B (Multiplier[12]));
XNOR2_X1 slo__sro_c356 (.ZN (p_1[12]), .A (slo__sro_n496), .B (n_12));
NAND2_X1 slo__sro_c375 (.ZN (slo__sro_n539), .A1 (Multiplier[21]), .A2 (n_21));
OAI21_X1 slo__sro_c376 (.ZN (slo__sro_n538), .A (p_0[21]), .B1 (n_21), .B2 (Multiplier[21]));
NAND2_X1 slo__sro_c377 (.ZN (n_22), .A1 (slo__sro_n539), .A2 (slo__sro_n538));
XNOR2_X1 slo__sro_c378 (.ZN (slo__sro_n537), .A (n_21), .B (Multiplier[21]));
XNOR2_X1 slo__sro_c379 (.ZN (p_1[21]), .A (slo__sro_n537), .B (p_0[21]));
NAND2_X1 slo__sro_c549 (.ZN (slo__sro_n755), .A1 (p_0[16]), .A2 (Multiplier[16]));
NOR2_X1 CLOCK_slo__sro_c977 (.ZN (CLOCK_slo__sro_n1567), .A1 (p_0[28]), .A2 (Multiplier[28]));
OAI21_X2 slo__sro_c551 (.ZN (n_17), .A (slo__sro_n755), .B1 (slo__sro_n756), .B2 (slo__sro_n754));
XNOR2_X2 slo__sro_c552 (.ZN (slo__sro_n753), .A (p_0[16]), .B (Multiplier[16]));
XNOR2_X1 slo__sro_c553 (.ZN (p_1[16]), .A (n_16), .B (slo__sro_n753));
NAND2_X1 CLOCK_slo__sro_c976 (.ZN (CLOCK_slo__sro_n1568), .A1 (p_0[28]), .A2 (Multiplier[28]));
OAI21_X1 CLOCK_slo__sro_c978 (.ZN (CLOCK_slo__sro_n1566), .A (CLOCK_slo__sro_n1568)
    , .B1 (CLOCK_slo__sro_n1567), .B2 (CLOCK_slo__sro_n1569));
XNOR2_X2 CLOCK_slo__sro_c979 (.ZN (CLOCK_slo__sro_n1565), .A (p_0[28]), .B (Multiplier[28]));
XNOR2_X1 CLOCK_slo__sro_c980 (.ZN (p_1[28]), .A (CLOCK_slo__sro_n1565), .B (n_28));
XNOR2_X2 CLOCK_slo__mro_c992 (.ZN (p_1[22]), .A (CLOCK_slo__mro_n1584), .B (p_0[22]));
NOR2_X1 CLOCK_slo__sro_c1003 (.ZN (CLOCK_slo__sro_n1598), .A1 (p_0[27]), .A2 (Multiplier[27]));
OAI21_X1 CLOCK_slo__sro_c1004 (.ZN (n_28), .A (CLOCK_slo__sro_n1599), .B1 (CLOCK_slo__sro_n1598), .B2 (CLOCK_slo__sro_n1600));
XNOR2_X1 CLOCK_slo__sro_c1005 (.ZN (CLOCK_slo__sro_n1597), .A (p_0[27]), .B (Multiplier[27]));
XNOR2_X1 CLOCK_slo__sro_c1006 (.ZN (p_1[27]), .A (CLOCK_slo__sro_n1597), .B (CLOCK_slo__sro_n1683));
INV_X1 CLOCK_slo__sro_c1022 (.ZN (CLOCK_slo__sro_n1622), .A (p_0[30]));
INV_X1 CLOCK_slo__sro_c1023 (.ZN (CLOCK_slo__sro_n1621), .A (n_30));
NOR2_X1 CLOCK_slo__sro_c1024 (.ZN (CLOCK_slo__sro_n1620), .A1 (n_33), .A2 (Multiplier[30]));
NAND2_X1 CLOCK_slo__sro_c1025 (.ZN (CLOCK_slo__sro_n1619), .A1 (CLOCK_slo__sro_n1621), .A2 (CLOCK_slo__sro_n1620));
NAND2_X1 CLOCK_slo__sro_c1026 (.ZN (CLOCK_slo__sro_n1618), .A1 (CLOCK_slo__sro_n1622), .A2 (CLOCK_slo__sro_n1623));
OAI21_X1 CLOCK_slo__sro_c1027 (.ZN (n_31), .A (CLOCK_slo__sro_n1619), .B1 (n_32), .B2 (CLOCK_slo__sro_n1618));
OAI21_X1 CLOCK_slo__sro_c1103 (.ZN (CLOCK_slo__sro_n1684), .A (p_0[26]), .B1 (CLOCK_slo__sro_n1860), .B2 (Multiplier[26]));
NAND2_X1 CLOCK_slo__sro_c1104 (.ZN (CLOCK_slo__sro_n1683), .A1 (CLOCK_slo__sro_n1684), .A2 (CLOCK_slo__sro_n1685));
XNOR2_X1 CLOCK_slo__sro_c1105 (.ZN (CLOCK_slo__sro_n1682), .A (CLOCK_slo__sro_n1860), .B (Multiplier[26]));
INV_X1 CLOCK_slo__xsl_c1067 (.ZN (CLOCK_slo__xsl_n1652), .A (n_9));
AND3_X4 CLOCK_slo__xsl_c1070 (.ZN (n_9), .A1 (slo__sro_n280), .A2 (slo__sro_n281), .A3 (slo__sro_n282));
INV_X1 CLOCK_slo__mro_c1143 (.ZN (CLOCK_slo__mro_n1722), .A (CLOCK_slo__mro_n1723));
XNOR2_X2 CLOCK_slo__mro_c1144 (.ZN (CLOCK_slo__mro_n1721), .A (p_0[8]), .B (slo__mro_n1013));
XNOR2_X1 CLOCK_slo__mro_c1145 (.ZN (p_1[8]), .A (CLOCK_slo__mro_n1721), .B (CLOCK_slo__mro_n1722));
XNOR2_X1 CLOCK_slo__sro_c1213 (.ZN (p_1[20]), .A (slo__sro_n245), .B (p_0[20]));
OAI21_X2 CLOCK_slo__sro_c1341 (.ZN (n_24), .A (slo__sro_n76), .B1 (slo__sro_n75), .B2 (slo__sro_n77));
OAI21_X2 CLOCK_slo__sro_c1255 (.ZN (CLOCK_slo__sro_n1860), .A (slo__sro_n200), .B1 (slo__sro_n199), .B2 (slo__sro_n201));

endmodule //datapath__0_176

module datapath__0_172 (p_0, p_1, p_2);

output [31:0] p_2;
input [31:0] p_0;
input [31:0] p_1;
wire slo__sro_n674;
wire CLOCK_slo__sro_n910;
wire n_1;
wire n_2;
wire n_3;
wire n_4;
wire n_7;
wire n_8;
wire n_9;
wire n_10;
wire n_11;
wire n_12;
wire n_13;
wire n_15;
wire n_17;
wire n_19;
wire n_20;
wire n_21;
wire n_22;
wire n_24;
wire n_26;
wire n_27;
wire n_28;
wire n_29;
wire n_30;
wire n_32;
wire n_0;
wire n_34;
wire n_33;
wire n_31;
wire slo__sro_n67;
wire slo__sro_n68;
wire slo__sro_n69;
wire slo__sro_n70;
wire slo__sro_n71;
wire slo__sro_n139;
wire slo__sro_n140;
wire slo__sro_n141;
wire slo__sro_n142;
wire slo__sro_n96;
wire slo__sro_n97;
wire slo__sro_n98;
wire slo__sro_n99;
wire slo__sro_n143;
wire slo__sro_n231;
wire slo__sro_n232;
wire slo__sro_n233;
wire slo__sro_n234;
wire slo__sro_n169;
wire slo__sro_n170;
wire slo__sro_n171;
wire slo__sro_n172;
wire slo__sro_n173;
wire slo__sro_n274;
wire slo__sro_n275;
wire slo__sro_n276;
wire slo__sro_n277;
wire slo__sro_n289;
wire slo__sro_n290;
wire slo__sro_n291;
wire slo__sro_n292;
wire slo__sro_n477;
wire slo__sro_n478;
wire slo__sro_n479;
wire slo__sro_n480;
wire slo__sro_n481;
wire slo__sro_n375;
wire slo__sro_n376;
wire slo__sro_n377;
wire slo__sro_n378;
wire slo__sro_n675;
wire slo__sro_n676;
wire slo__sro_n677;
wire CLOCK_slo__sro_n911;
wire CLOCK_slo__sro_n912;
wire CLOCK_slo__sro_n913;
wire CLOCK_slo__sro_n914;
wire CLOCK_slo__sro_n915;
wire CLOCK_slo__sro_n1177;
wire CLOCK_slo__sro_n1178;
wire CLOCK_slo__sro_n1179;
wire CLOCK_slo__sro_n1180;
wire CLOCK_slo__sro_n1080;
wire CLOCK_slo__sro_n1081;
wire CLOCK_slo__sro_n1082;
wire CLOCK_slo__sro_n1083;
wire CLOCK_slo__sro_n979;
wire CLOCK_slo__sro_n980;
wire CLOCK_slo__sro_n981;
wire CLOCK_slo__sro_n982;
wire CLOCK_slo__sro_n1200;
wire CLOCK_slo__sro_n1745;
wire CLOCK_slo__sro_n1746;
wire CLOCK_slo__sro_n1747;
wire CLOCK_slo__sro_n1748;
wire CLOCK_slo__sro_n1749;
wire CLOCK_slo__sro_n1619;
wire CLOCK_slo__sro_n1620;
wire CLOCK_slo__sro_n1621;
wire CLOCK_slo__sro_n1622;


INV_X1 i_36 (.ZN (n_34), .A (p_0[30]));
INV_X1 i_35 (.ZN (n_33), .A (p_1[30]));
INV_X1 i_34 (.ZN (n_32), .A (n_30));
XOR2_X1 i_32 (.Z (p_2[31]), .A (p_0[31]), .B (n_31));
OAI22_X1 i_31 (.ZN (n_0), .A1 (n_34), .A2 (p_1[30]), .B1 (p_0[30]), .B2 (n_33));
XNOR2_X1 i_0 (.ZN (p_2[30]), .A (n_32), .B (n_0));
FA_X1 i_30 (.CO (n_30), .S (p_2[29]), .A (p_0[29]), .B (p_1[29]), .CI (n_29));
FA_X1 i_28 (.CO (n_28), .S (p_2[27]), .A (p_0[27]), .B (p_1[27]), .CI (n_27));
FA_X1 i_27 (.CO (n_27), .S (p_2[26]), .A (p_0[26]), .B (p_1[26]), .CI (n_26));
FA_X1 i_26 (.CO (n_26), .S (p_2[25]), .A (p_0[25]), .B (p_1[25]), .CI (slo__sro_n68));
INV_X1 slo__sro_c72 (.ZN (slo__sro_n143), .A (n_22));
FA_X1 i_24 (.CO (n_24), .S (p_2[23]), .A (p_0[23]), .B (p_1[23]), .CI (slo__sro_n140));
INV_X1 slo__sro_c152 (.ZN (slo__sro_n234), .A (CLOCK_slo__sro_n1746));
FA_X1 i_22 (.CO (n_22), .S (p_2[21]), .A (p_0[21]), .B (p_1[21]), .CI (n_21));
FA_X1 i_20 (.CO (n_20), .S (p_2[19]), .A (p_0[19]), .B (p_1[19]), .CI (n_19));
INV_X2 slo__sro_c194 (.ZN (slo__sro_n277), .A (n_11));
NAND2_X1 slo__sro_c153 (.ZN (slo__sro_n233), .A1 (p_1[18]), .A2 (p_0[18]));
NAND2_X1 slo__sro_c423 (.ZN (slo__sro_n675), .A1 (slo__sro_n676), .A2 (slo__sro_n677));
FA_X1 i_15 (.CO (n_15), .S (p_2[14]), .A (p_0[14]), .B (p_1[14]), .CI (slo__sro_n478));
NAND2_X1 slo__sro_c421 (.ZN (slo__sro_n677), .A1 (slo__sro_n170), .A2 (p_0[5]));
FA_X1 i_13 (.CO (n_13), .S (p_2[12]), .A (p_0[12]), .B (p_1[12]), .CI (n_12));
INV_X1 slo__sro_c208 (.ZN (slo__sro_n292), .A (n_7));
FA_X1 i_10 (.CO (n_10), .S (p_2[9]), .A (p_0[9]), .B (p_1[9]), .CI (n_9));
INV_X1 slo__sro_c339 (.ZN (slo__sro_n481), .A (p_1[13]));
FA_X1 i_7 (.CO (n_7), .S (p_2[6]), .A (p_0[6]), .B (p_1[6]), .CI (slo__sro_n675));
INV_X1 CLOCK_slo__sro_c533 (.ZN (CLOCK_slo__sro_n915), .A (n_34));
NAND2_X1 slo__sro_c195 (.ZN (slo__sro_n276), .A1 (p_1[11]), .A2 (p_0[11]));
FA_X1 i_4 (.CO (n_4), .S (p_2[3]), .A (p_0[3]), .B (p_1[3]), .CI (n_3));
FA_X1 i_3 (.CO (n_3), .S (p_2[2]), .A (p_0[2]), .B (p_1[2]), .CI (n_2));
FA_X1 i_2 (.CO (n_2), .S (p_2[1]), .A (p_0[1]), .B (p_1[1]), .CI (n_1));
HA_X1 i_1 (.CO (n_1), .S (p_2[0]), .A (p_0[0]), .B (p_1[0]));
INV_X1 slo__sro_c5 (.ZN (slo__sro_n71), .A (n_24));
NAND2_X1 slo__sro_c6 (.ZN (slo__sro_n70), .A1 (p_1[24]), .A2 (p_0[24]));
NOR2_X1 slo__sro_c7 (.ZN (slo__sro_n69), .A1 (p_1[24]), .A2 (p_0[24]));
OAI21_X1 slo__sro_c8 (.ZN (slo__sro_n68), .A (slo__sro_n70), .B1 (slo__sro_n71), .B2 (slo__sro_n69));
XNOR2_X1 slo__sro_c9 (.ZN (slo__sro_n67), .A (p_1[24]), .B (p_0[24]));
XNOR2_X1 slo__sro_c10 (.ZN (p_2[24]), .A (slo__sro_n67), .B (n_24));
NAND2_X1 slo__sro_c73 (.ZN (slo__sro_n142), .A1 (p_1[22]), .A2 (p_0[22]));
NOR2_X1 slo__sro_c74 (.ZN (slo__sro_n141), .A1 (p_1[22]), .A2 (p_0[22]));
OAI21_X1 slo__sro_c75 (.ZN (slo__sro_n140), .A (slo__sro_n142), .B1 (slo__sro_n143), .B2 (slo__sro_n141));
XNOR2_X1 slo__sro_c76 (.ZN (slo__sro_n139), .A (p_1[22]), .B (p_0[22]));
XNOR2_X1 slo__sro_c77 (.ZN (p_2[22]), .A (slo__sro_n139), .B (n_22));
INV_X1 slo__sro_c32 (.ZN (slo__sro_n99), .A (CLOCK_slo__sro_n1200));
NAND2_X1 slo__sro_c33 (.ZN (slo__sro_n98), .A1 (p_1[16]), .A2 (p_0[16]));
NOR2_X1 slo__sro_c34 (.ZN (slo__sro_n97), .A1 (p_1[16]), .A2 (p_0[16]));
OAI21_X1 slo__sro_c35 (.ZN (n_17), .A (slo__sro_n98), .B1 (slo__sro_n99), .B2 (slo__sro_n97));
XNOR2_X1 slo__sro_c36 (.ZN (slo__sro_n96), .A (p_1[16]), .B (p_0[16]));
XNOR2_X1 slo__sro_c37 (.ZN (p_2[16]), .A (slo__sro_n96), .B (CLOCK_slo__sro_n1200));
NOR2_X1 slo__sro_c154 (.ZN (slo__sro_n232), .A1 (p_1[18]), .A2 (p_0[18]));
OAI21_X1 slo__sro_c155 (.ZN (n_19), .A (slo__sro_n233), .B1 (slo__sro_n234), .B2 (slo__sro_n232));
XNOR2_X1 slo__sro_c156 (.ZN (slo__sro_n231), .A (p_1[18]), .B (p_0[18]));
XNOR2_X1 slo__sro_c157 (.ZN (p_2[18]), .A (slo__sro_n231), .B (CLOCK_slo__sro_n1746));
INV_X1 slo__sro_c99 (.ZN (slo__sro_n173), .A (n_4));
NAND2_X1 slo__sro_c100 (.ZN (slo__sro_n172), .A1 (p_1[4]), .A2 (p_0[4]));
NOR2_X1 slo__sro_c101 (.ZN (slo__sro_n171), .A1 (p_1[4]), .A2 (p_0[4]));
OAI21_X2 slo__sro_c102 (.ZN (slo__sro_n170), .A (slo__sro_n172), .B1 (slo__sro_n171), .B2 (slo__sro_n173));
XNOR2_X2 slo__sro_c103 (.ZN (slo__sro_n169), .A (p_1[4]), .B (p_0[4]));
XNOR2_X2 slo__sro_c104 (.ZN (p_2[4]), .A (slo__sro_n169), .B (n_4));
NOR2_X1 slo__sro_c196 (.ZN (slo__sro_n275), .A1 (p_1[11]), .A2 (p_0[11]));
OAI21_X2 slo__sro_c197 (.ZN (n_12), .A (slo__sro_n276), .B1 (slo__sro_n277), .B2 (slo__sro_n275));
XNOR2_X1 slo__sro_c198 (.ZN (slo__sro_n274), .A (p_1[11]), .B (p_0[11]));
NAND2_X1 slo__sro_c209 (.ZN (slo__sro_n291), .A1 (p_1[7]), .A2 (p_0[7]));
NOR2_X1 slo__sro_c210 (.ZN (slo__sro_n290), .A1 (p_1[7]), .A2 (p_0[7]));
OAI21_X1 slo__sro_c211 (.ZN (n_8), .A (slo__sro_n291), .B1 (slo__sro_n292), .B2 (slo__sro_n290));
XNOR2_X2 slo__sro_c212 (.ZN (slo__sro_n289), .A (p_1[7]), .B (p_0[7]));
XNOR2_X2 slo__sro_c213 (.ZN (p_2[7]), .A (slo__sro_n289), .B (n_7));
NAND2_X1 slo__sro_c340 (.ZN (slo__sro_n480), .A1 (n_13), .A2 (p_0[13]));
NOR2_X2 slo__sro_c341 (.ZN (slo__sro_n479), .A1 (n_13), .A2 (p_0[13]));
OAI21_X1 slo__sro_c342 (.ZN (slo__sro_n478), .A (slo__sro_n480), .B1 (slo__sro_n479), .B2 (slo__sro_n481));
XNOR2_X1 slo__sro_c343 (.ZN (slo__sro_n477), .A (n_13), .B (p_0[13]));
XNOR2_X1 slo__sro_c344 (.ZN (p_2[13]), .A (slo__sro_n477), .B (p_1[13]));
OAI21_X1 slo__sro_c422 (.ZN (slo__sro_n676), .A (p_1[5]), .B1 (slo__sro_n170), .B2 (p_0[5]));
INV_X1 slo__sro_c255 (.ZN (slo__sro_n378), .A (n_15));
NAND2_X1 slo__sro_c256 (.ZN (slo__sro_n377), .A1 (p_1[15]), .A2 (p_0[15]));
NOR2_X1 slo__sro_c257 (.ZN (slo__sro_n376), .A1 (p_1[15]), .A2 (p_0[15]));
XNOR2_X1 slo__sro_c259 (.ZN (slo__sro_n375), .A (p_1[15]), .B (p_0[15]));
XNOR2_X1 slo__sro_c260 (.ZN (p_2[15]), .A (slo__sro_n375), .B (n_15));
XNOR2_X2 slo__sro_c424 (.ZN (slo__sro_n674), .A (slo__sro_n170), .B (p_0[5]));
XNOR2_X1 slo__sro_c425 (.ZN (p_2[5]), .A (slo__sro_n674), .B (p_1[5]));
INV_X1 CLOCK_slo__sro_c534 (.ZN (CLOCK_slo__sro_n914), .A (p_1[30]));
INV_X1 CLOCK_slo__sro_c535 (.ZN (CLOCK_slo__sro_n913), .A (n_30));
NOR2_X1 CLOCK_slo__sro_c536 (.ZN (CLOCK_slo__sro_n912), .A1 (n_33), .A2 (p_0[30]));
NAND2_X1 CLOCK_slo__sro_c537 (.ZN (CLOCK_slo__sro_n911), .A1 (CLOCK_slo__sro_n913), .A2 (CLOCK_slo__sro_n912));
NAND2_X1 CLOCK_slo__sro_c538 (.ZN (CLOCK_slo__sro_n910), .A1 (CLOCK_slo__sro_n914), .A2 (CLOCK_slo__sro_n915));
OAI21_X1 CLOCK_slo__sro_c539 (.ZN (n_31), .A (CLOCK_slo__sro_n911), .B1 (n_32), .B2 (CLOCK_slo__sro_n910));
INV_X1 CLOCK_slo__sro_c827 (.ZN (CLOCK_slo__sro_n1180), .A (n_8));
NAND2_X1 CLOCK_slo__sro_c828 (.ZN (CLOCK_slo__sro_n1179), .A1 (p_1[8]), .A2 (p_0[8]));
NOR2_X1 CLOCK_slo__sro_c829 (.ZN (CLOCK_slo__sro_n1178), .A1 (p_1[8]), .A2 (p_0[8]));
OAI21_X1 CLOCK_slo__sro_c830 (.ZN (n_9), .A (CLOCK_slo__sro_n1179), .B1 (CLOCK_slo__sro_n1180), .B2 (CLOCK_slo__sro_n1178));
XNOR2_X1 CLOCK_slo__sro_c831 (.ZN (CLOCK_slo__sro_n1177), .A (p_1[8]), .B (p_0[8]));
XNOR2_X1 CLOCK_slo__sro_c832 (.ZN (p_2[8]), .A (CLOCK_slo__sro_n1177), .B (n_8));
INV_X1 CLOCK_slo__sro_c727 (.ZN (CLOCK_slo__sro_n1083), .A (n_28));
NAND2_X1 CLOCK_slo__sro_c728 (.ZN (CLOCK_slo__sro_n1082), .A1 (p_1[28]), .A2 (p_0[28]));
NOR2_X1 CLOCK_slo__sro_c729 (.ZN (CLOCK_slo__sro_n1081), .A1 (p_1[28]), .A2 (p_0[28]));
OAI21_X1 CLOCK_slo__sro_c730 (.ZN (n_29), .A (CLOCK_slo__sro_n1082), .B1 (CLOCK_slo__sro_n1083), .B2 (CLOCK_slo__sro_n1081));
XNOR2_X1 CLOCK_slo__sro_c731 (.ZN (CLOCK_slo__sro_n1080), .A (p_1[28]), .B (p_0[28]));
XNOR2_X1 CLOCK_slo__sro_c732 (.ZN (p_2[28]), .A (CLOCK_slo__sro_n1080), .B (n_28));
OAI21_X1 CLOCK_slo__sro_c851 (.ZN (CLOCK_slo__sro_n1200), .A (slo__sro_n377), .B1 (slo__sro_n378), .B2 (slo__sro_n376));
XNOR2_X1 CLOCK_slo__sro_c983 (.ZN (p_2[11]), .A (n_11), .B (slo__sro_n274));
INV_X2 CLOCK_slo__sro_c624 (.ZN (CLOCK_slo__sro_n982), .A (n_10));
NAND2_X1 CLOCK_slo__sro_c625 (.ZN (CLOCK_slo__sro_n981), .A1 (p_1[10]), .A2 (p_0[10]));
NOR2_X1 CLOCK_slo__sro_c626 (.ZN (CLOCK_slo__sro_n980), .A1 (p_1[10]), .A2 (p_0[10]));
OAI21_X2 CLOCK_slo__sro_c627 (.ZN (n_11), .A (CLOCK_slo__sro_n981), .B1 (CLOCK_slo__sro_n982), .B2 (CLOCK_slo__sro_n980));
XNOR2_X1 CLOCK_slo__sro_c628 (.ZN (CLOCK_slo__sro_n979), .A (p_1[10]), .B (p_0[10]));
XNOR2_X1 CLOCK_slo__sro_c629 (.ZN (p_2[10]), .A (CLOCK_slo__sro_n979), .B (n_10));
INV_X1 CLOCK_slo__sro_c1433 (.ZN (CLOCK_slo__sro_n1749), .A (n_17));
NAND2_X1 CLOCK_slo__sro_c1434 (.ZN (CLOCK_slo__sro_n1748), .A1 (p_1[17]), .A2 (p_0[17]));
NOR2_X1 CLOCK_slo__sro_c1435 (.ZN (CLOCK_slo__sro_n1747), .A1 (p_1[17]), .A2 (p_0[17]));
OAI21_X1 CLOCK_slo__sro_c1436 (.ZN (CLOCK_slo__sro_n1746), .A (CLOCK_slo__sro_n1748)
    , .B1 (CLOCK_slo__sro_n1749), .B2 (CLOCK_slo__sro_n1747));
XNOR2_X2 CLOCK_slo__sro_c1437 (.ZN (CLOCK_slo__sro_n1745), .A (p_1[17]), .B (p_0[17]));
XNOR2_X1 CLOCK_slo__sro_c1438 (.ZN (p_2[17]), .A (CLOCK_slo__sro_n1745), .B (n_17));
INV_X1 CLOCK_slo__sro_c1284 (.ZN (CLOCK_slo__sro_n1622), .A (n_20));
NAND2_X1 CLOCK_slo__sro_c1285 (.ZN (CLOCK_slo__sro_n1621), .A1 (p_1[20]), .A2 (p_0[20]));
NOR2_X1 CLOCK_slo__sro_c1286 (.ZN (CLOCK_slo__sro_n1620), .A1 (p_1[20]), .A2 (p_0[20]));
OAI21_X1 CLOCK_slo__sro_c1287 (.ZN (n_21), .A (CLOCK_slo__sro_n1621), .B1 (CLOCK_slo__sro_n1622), .B2 (CLOCK_slo__sro_n1620));
XNOR2_X1 CLOCK_slo__sro_c1288 (.ZN (CLOCK_slo__sro_n1619), .A (p_1[20]), .B (p_0[20]));
XNOR2_X1 CLOCK_slo__sro_c1289 (.ZN (p_2[20]), .A (CLOCK_slo__sro_n1619), .B (n_20));

endmodule //datapath__0_172

module datapath__0_171 (Multiplier, p_0, p_1);

output [31:0] p_1;
input [31:0] Multiplier;
input [31:0] p_0;
wire CLOCK_slo__mro_n1682;
wire n_1;
wire n_2;
wire n_3;
wire n_4;
wire n_5;
wire n_6;
wire n_7;
wire n_8;
wire n_9;
wire n_11;
wire CLOCK_slo__mro_n1258;
wire n_14;
wire n_15;
wire n_17;
wire n_18;
wire n_19;
wire n_20;
wire CLOCK_slo__sro_n1359;
wire n_22;
wire n_23;
wire n_25;
wire n_27;
wire n_28;
wire n_30;
wire n_32;
wire n_0;
wire n_34;
wire n_33;
wire n_31;
wire slo__sro_n59;
wire slo__sro_n60;
wire slo__sro_n61;
wire slo__sro_n62;
wire slo__sro_n63;
wire slo__sro_n77;
wire slo__sro_n78;
wire slo__sro_n79;
wire slo__sro_n89;
wire slo__sro_n90;
wire slo__sro_n91;
wire slo__sro_n92;
wire slo__sro_n105;
wire slo__sro_n106;
wire slo__sro_n115;
wire slo__sro_n116;
wire slo__sro_n117;
wire slo__sro_n118;
wire slo__sro_n119;
wire slo__sro_n132;
wire slo__sro_n133;
wire slo__sro_n134;
wire slo__sro_n135;
wire CLOCK_slo__sro_n1465;
wire slo__sro_n162;
wire slo__sro_n163;
wire slo__sro_n164;
wire slo__sro_n193;
wire slo__sro_n194;
wire slo__sro_n195;
wire slo__sro_n196;
wire slo__sro_n197;
wire slo__sro_n210;
wire slo__sro_n211;
wire slo__sro_n212;
wire slo__sro_n213;
wire slo__sro_n229;
wire slo__sro_n230;
wire slo__sro_n231;
wire slo__sro_n232;
wire slo__sro_n247;
wire slo__sro_n248;
wire slo__mro_n698;
wire slo__mro_n699;
wire slo__mro_n756;
wire slo__mro_n700;
wire slo__mro_n701;
wire CLOCK_slo__sro_n1360;
wire CLOCK_slo__sro_n1361;
wire CLOCK_slo__sro_n1362;
wire CLOCK_slo__sro_n1389;
wire CLOCK_slo__sro_n1390;
wire CLOCK_slo__sro_n1391;
wire CLOCK_slo__sro_n1392;
wire CLOCK_slo__sro_n1393;
wire CLOCK_slo__sro_n1408;
wire CLOCK_slo__sro_n1409;
wire CLOCK_slo__sro_n1410;
wire CLOCK_slo__sro_n1411;
wire CLOCK_slo__xsl_n1441;
wire CLOCK_slo__sro_n1466;
wire slo__sro_n831;
wire slo__sro_n832;
wire slo__sro_n833;
wire slo__sro_n834;
wire CLOCK_slo__sro_n1467;
wire CLOCK_slo__sro_n1468;
wire CLOCK_slo__sro_n1493;
wire CLOCK_slo__sro_n1494;
wire CLOCK_slo__sro_n1495;
wire CLOCK_slo__sro_n1496;
wire CLOCK_slo__sro_n1660;
wire CLOCK_slo__sro_n1661;
wire CLOCK_slo__xsl_n1561;
wire CLOCK_slo__xsl_n1562;
wire CLOCK_slo__sro_n1613;
wire CLOCK_slo__sro_n1614;
wire CLOCK_slo__sro_n1615;
wire CLOCK_slo__sro_n1616;


INV_X1 i_36 (.ZN (n_34), .A (Multiplier[30]));
INV_X1 i_35 (.ZN (n_33), .A (p_0[30]));
INV_X1 i_34 (.ZN (n_32), .A (n_30));
XOR2_X1 i_32 (.Z (p_1[31]), .A (Multiplier[31]), .B (n_31));
OAI22_X1 i_31 (.ZN (n_0), .A1 (n_34), .A2 (p_0[30]), .B1 (Multiplier[30]), .B2 (n_33));
XNOR2_X1 i_0 (.ZN (p_1[30]), .A (n_32), .B (n_0));
FA_X1 i_30 (.CO (n_30), .S (p_1[29]), .A (Multiplier[29]), .B (p_0[29]), .CI (CLOCK_slo__sro_n1360));
INV_X1 CLOCK_slo__sro_c1005 (.ZN (CLOCK_slo__sro_n1393), .A (n_23));
FA_X1 i_28 (.CO (n_28), .S (p_1[27]), .A (Multiplier[27]), .B (p_0[27]), .CI (n_27));
FA_X1 i_27 (.CO (n_27), .S (p_1[26]), .A (Multiplier[26]), .B (p_0[26]), .CI (slo__sro_n162));
INV_X1 slo__sro_c123 (.ZN (slo__sro_n197), .A (n_15));
INV_X1 slo__sro_c29 (.ZN (slo__sro_n92), .A (slo__sro_n194));
INV_X1 CLOCK_slo__sro_c1021 (.ZN (CLOCK_slo__sro_n1411), .A (n_17));
FA_X1 i_23 (.CO (n_23), .S (p_1[22]), .A (Multiplier[22]), .B (p_0[22]), .CI (n_22));
INV_X1 slo__sro_c55 (.ZN (slo__sro_n119), .A (n_9));
INV_X1 slo__sro_c15 (.ZN (slo__sro_n79), .A (CLOCK_slo__sro_n1390));
FA_X1 i_20 (.CO (n_20), .S (p_1[19]), .A (Multiplier[19]), .B (p_0[19]), .CI (n_19));
NAND2_X1 CLOCK_slo__sro_c1128 (.ZN (CLOCK_slo__sro_n1495), .A1 (n_5), .A2 (Multiplier[5]));
INV_X1 CLOCK_slo__sro_c1100 (.ZN (CLOCK_slo__sro_n1468), .A (n_3));
NAND2_X1 slo__sro_c43 (.ZN (slo__sro_n106), .A1 (slo__sro_n60), .A2 (Multiplier[21]));
NAND2_X1 slo__sro_c137 (.ZN (slo__sro_n213), .A1 (p_0[13]), .A2 (Multiplier[13]));
FA_X1 i_15 (.CO (n_15), .S (p_1[14]), .A (Multiplier[14]), .B (p_0[14]), .CI (n_14));
INV_X1 slo__sro_c155 (.ZN (slo__sro_n232), .A (n_8));
NAND2_X1 slo__sro_c96 (.ZN (slo__sro_n164), .A1 (n_25), .A2 (Multiplier[25]));
INV_X1 slo__mro_c499 (.ZN (slo__mro_n701), .A (Multiplier[25]));
NOR2_X1 CLOCK_slo__sro_c1102 (.ZN (CLOCK_slo__sro_n1466), .A1 (p_0[3]), .A2 (Multiplier[3]));
NAND2_X1 slo__sro_c171 (.ZN (slo__sro_n248), .A1 (slo__sro_n116), .A2 (Multiplier[10]));
FA_X1 i_8 (.CO (n_8), .S (p_1[7]), .A (Multiplier[7]), .B (p_0[7]), .CI (n_7));
FA_X1 i_7 (.CO (n_7), .S (p_1[6]), .A (Multiplier[6]), .B (p_0[6]), .CI (n_6));
OR2_X1 CLOCK_slo__sro_c1282 (.ZN (CLOCK_slo__sro_n1661), .A1 (n_33), .A2 (Multiplier[30]));
FA_X1 i_5 (.CO (n_5), .S (p_1[4]), .A (Multiplier[4]), .B (p_0[4]), .CI (n_4));
INV_X1 CLOCK_slo__sro_c1127 (.ZN (CLOCK_slo__sro_n1496), .A (p_0[5]));
FA_X1 i_3 (.CO (n_3), .S (p_1[2]), .A (Multiplier[2]), .B (p_0[2]), .CI (n_2));
FA_X1 i_2 (.CO (n_2), .S (p_1[1]), .A (Multiplier[1]), .B (p_0[1]), .CI (n_1));
HA_X1 i_1 (.CO (n_1), .S (p_1[0]), .A (Multiplier[0]), .B (p_0[0]));
INV_X1 slo__sro_c1 (.ZN (slo__sro_n63), .A (n_20));
NAND2_X1 slo__sro_c2 (.ZN (slo__sro_n62), .A1 (p_0[20]), .A2 (Multiplier[20]));
NOR2_X1 slo__sro_c3 (.ZN (slo__sro_n61), .A1 (p_0[20]), .A2 (Multiplier[20]));
OAI21_X1 slo__sro_c4 (.ZN (slo__sro_n60), .A (slo__sro_n62), .B1 (slo__sro_n63), .B2 (slo__sro_n61));
XNOR2_X1 slo__sro_c5 (.ZN (slo__sro_n59), .A (p_0[20]), .B (Multiplier[20]));
XNOR2_X2 slo__sro_c6 (.ZN (p_1[20]), .A (slo__sro_n59), .B (n_20));
NAND2_X1 slo__sro_c16 (.ZN (slo__sro_n78), .A1 (p_0[24]), .A2 (Multiplier[24]));
NOR2_X1 slo__sro_c17 (.ZN (slo__sro_n77), .A1 (p_0[24]), .A2 (Multiplier[24]));
OAI21_X1 slo__sro_c18 (.ZN (n_25), .A (slo__sro_n78), .B1 (slo__sro_n79), .B2 (slo__sro_n77));
NAND2_X1 CLOCK_slo__sro_c980 (.ZN (CLOCK_slo__sro_n1362), .A1 (p_0[28]), .A2 (Multiplier[28]));
OAI21_X1 CLOCK_slo__sro_c981 (.ZN (CLOCK_slo__sro_n1361), .A (n_28), .B1 (p_0[28]), .B2 (Multiplier[28]));
NAND2_X1 slo__sro_c30 (.ZN (slo__sro_n91), .A1 (p_0[16]), .A2 (Multiplier[16]));
NOR2_X1 slo__sro_c31 (.ZN (slo__sro_n90), .A1 (p_0[16]), .A2 (Multiplier[16]));
OAI21_X1 slo__sro_c32 (.ZN (n_17), .A (slo__sro_n91), .B1 (slo__sro_n92), .B2 (slo__sro_n90));
XNOR2_X1 slo__sro_c33 (.ZN (slo__sro_n89), .A (p_0[16]), .B (Multiplier[16]));
XNOR2_X2 slo__sro_c34 (.ZN (p_1[16]), .A (slo__sro_n89), .B (slo__sro_n194));
OAI21_X1 slo__sro_c44 (.ZN (slo__sro_n105), .A (p_0[21]), .B1 (slo__sro_n60), .B2 (Multiplier[21]));
NAND2_X1 slo__sro_c45 (.ZN (n_22), .A1 (slo__sro_n105), .A2 (slo__sro_n106));
XNOR2_X1 CLOCK_slo__mro_c1316 (.ZN (p_1[10]), .A (CLOCK_slo__mro_n1682), .B (slo__sro_n116));
XNOR2_X1 CLOCK_slo__mro_c1315 (.ZN (CLOCK_slo__mro_n1682), .A (p_0[10]), .B (Multiplier[10]));
NAND2_X1 slo__sro_c56 (.ZN (slo__sro_n118), .A1 (p_0[9]), .A2 (Multiplier[9]));
NOR2_X2 slo__sro_c57 (.ZN (slo__sro_n117), .A1 (p_0[9]), .A2 (Multiplier[9]));
OAI21_X2 slo__sro_c58 (.ZN (slo__sro_n116), .A (slo__sro_n118), .B1 (slo__sro_n119), .B2 (slo__sro_n117));
XNOR2_X2 slo__sro_c59 (.ZN (slo__sro_n115), .A (p_0[9]), .B (Multiplier[9]));
XNOR2_X2 slo__sro_c60 (.ZN (p_1[9]), .A (slo__sro_n115), .B (CLOCK_slo__xsl_n1561));
NAND2_X1 slo__sro_c70 (.ZN (slo__sro_n135), .A1 (p_0[11]), .A2 (Multiplier[11]));
NOR2_X1 slo__sro_c71 (.ZN (slo__sro_n134), .A1 (p_0[11]), .A2 (Multiplier[11]));
OAI21_X1 slo__sro_c72 (.ZN (slo__sro_n133), .A (slo__sro_n135), .B1 (n_11), .B2 (slo__sro_n134));
XNOR2_X2 slo__sro_c73 (.ZN (slo__sro_n132), .A (p_0[11]), .B (Multiplier[11]));
XNOR2_X2 slo__sro_c74 (.ZN (p_1[11]), .A (slo__sro_n132), .B (CLOCK_slo__xsl_n1441));
OAI21_X1 slo__sro_c97 (.ZN (slo__sro_n163), .A (p_0[25]), .B1 (n_25), .B2 (Multiplier[25]));
NAND2_X1 slo__sro_c98 (.ZN (slo__sro_n162), .A1 (slo__sro_n163), .A2 (slo__sro_n164));
XNOR2_X1 slo__mro_c532 (.ZN (p_1[21]), .A (slo__mro_n756), .B (slo__sro_n60));
XNOR2_X2 CLOCK_slo__mro_c881 (.ZN (CLOCK_slo__mro_n1258), .A (p_0[24]), .B (Multiplier[24]));
NAND2_X1 slo__sro_c124 (.ZN (slo__sro_n196), .A1 (p_0[15]), .A2 (Multiplier[15]));
NOR2_X1 slo__sro_c125 (.ZN (slo__sro_n195), .A1 (p_0[15]), .A2 (Multiplier[15]));
OAI21_X1 slo__sro_c126 (.ZN (slo__sro_n194), .A (slo__sro_n196), .B1 (slo__sro_n197), .B2 (slo__sro_n195));
XNOR2_X2 slo__sro_c127 (.ZN (slo__sro_n193), .A (p_0[15]), .B (Multiplier[15]));
XNOR2_X1 slo__sro_c128 (.ZN (p_1[15]), .A (slo__sro_n193), .B (n_15));
NAND2_X1 slo__sro_c138 (.ZN (slo__sro_n212), .A1 (CLOCK_slo__sro_n1614), .A2 (Multiplier[13]));
NAND2_X1 slo__sro_c139 (.ZN (slo__sro_n211), .A1 (CLOCK_slo__sro_n1614), .A2 (p_0[13]));
NAND3_X1 slo__sro_c140 (.ZN (n_14), .A1 (slo__sro_n212), .A2 (slo__sro_n211), .A3 (slo__sro_n213));
XNOR2_X1 slo__sro_c141 (.ZN (slo__sro_n210), .A (p_0[13]), .B (Multiplier[13]));
XNOR2_X1 slo__sro_c142 (.ZN (p_1[13]), .A (slo__sro_n210), .B (CLOCK_slo__sro_n1614));
NAND2_X1 slo__sro_c156 (.ZN (slo__sro_n231), .A1 (p_0[8]), .A2 (Multiplier[8]));
NOR2_X1 slo__sro_c157 (.ZN (slo__sro_n230), .A1 (p_0[8]), .A2 (Multiplier[8]));
OAI21_X1 slo__sro_c158 (.ZN (n_9), .A (slo__sro_n231), .B1 (slo__sro_n232), .B2 (slo__sro_n230));
XNOR2_X2 slo__sro_c159 (.ZN (slo__sro_n229), .A (p_0[8]), .B (Multiplier[8]));
XNOR2_X1 slo__sro_c160 (.ZN (p_1[8]), .A (n_8), .B (slo__sro_n229));
OAI21_X2 slo__sro_c172 (.ZN (slo__sro_n247), .A (p_0[10]), .B1 (slo__sro_n116), .B2 (Multiplier[10]));
XNOR2_X2 CLOCK_slo__sro_c1104 (.ZN (CLOCK_slo__sro_n1465), .A (p_0[3]), .B (Multiplier[3]));
OAI21_X1 slo__mro_c500 (.ZN (slo__mro_n700), .A (slo__sro_n78), .B1 (slo__sro_n79), .B2 (slo__sro_n77));
INV_X1 slo__mro_c501 (.ZN (slo__mro_n699), .A (slo__mro_n700));
XNOR2_X2 slo__mro_c531 (.ZN (slo__mro_n756), .A (p_0[21]), .B (Multiplier[21]));
XNOR2_X1 slo__mro_c502 (.ZN (slo__mro_n698), .A (p_0[25]), .B (slo__mro_n701));
XNOR2_X2 slo__mro_c503 (.ZN (p_1[25]), .A (slo__mro_n698), .B (slo__mro_n699));
XNOR2_X1 CLOCK_slo__mro_c882 (.ZN (p_1[24]), .A (CLOCK_slo__mro_n1258), .B (CLOCK_slo__sro_n1390));
NAND2_X1 CLOCK_slo__sro_c982 (.ZN (CLOCK_slo__sro_n1360), .A1 (CLOCK_slo__sro_n1361), .A2 (CLOCK_slo__sro_n1362));
XNOR2_X2 CLOCK_slo__sro_c983 (.ZN (CLOCK_slo__sro_n1359), .A (p_0[28]), .B (Multiplier[28]));
XNOR2_X1 CLOCK_slo__sro_c984 (.ZN (p_1[28]), .A (CLOCK_slo__sro_n1359), .B (n_28));
NAND2_X1 CLOCK_slo__sro_c1006 (.ZN (CLOCK_slo__sro_n1392), .A1 (p_0[23]), .A2 (Multiplier[23]));
NOR2_X1 CLOCK_slo__sro_c1007 (.ZN (CLOCK_slo__sro_n1391), .A1 (p_0[23]), .A2 (Multiplier[23]));
OAI21_X1 CLOCK_slo__sro_c1008 (.ZN (CLOCK_slo__sro_n1390), .A (CLOCK_slo__sro_n1392)
    , .B1 (CLOCK_slo__sro_n1393), .B2 (CLOCK_slo__sro_n1391));
XNOR2_X1 CLOCK_slo__sro_c1009 (.ZN (CLOCK_slo__sro_n1389), .A (p_0[23]), .B (Multiplier[23]));
XNOR2_X1 CLOCK_slo__sro_c1010 (.ZN (p_1[23]), .A (CLOCK_slo__sro_n1389), .B (n_23));
NAND2_X1 CLOCK_slo__sro_c1022 (.ZN (CLOCK_slo__sro_n1410), .A1 (p_0[17]), .A2 (Multiplier[17]));
NOR2_X1 CLOCK_slo__sro_c1023 (.ZN (CLOCK_slo__sro_n1409), .A1 (p_0[17]), .A2 (Multiplier[17]));
OAI21_X2 CLOCK_slo__sro_c1024 (.ZN (n_18), .A (CLOCK_slo__sro_n1410), .B1 (CLOCK_slo__sro_n1411), .B2 (CLOCK_slo__sro_n1409));
XNOR2_X1 CLOCK_slo__sro_c1025 (.ZN (CLOCK_slo__sro_n1408), .A (p_0[17]), .B (Multiplier[17]));
XNOR2_X1 CLOCK_slo__sro_c1026 (.ZN (p_1[17]), .A (CLOCK_slo__sro_n1408), .B (n_17));
NAND2_X1 CLOCK_slo__sro_c1101 (.ZN (CLOCK_slo__sro_n1467), .A1 (p_0[3]), .A2 (Multiplier[3]));
OAI21_X1 CLOCK_slo__sro_c1103 (.ZN (n_4), .A (CLOCK_slo__sro_n1467), .B1 (CLOCK_slo__sro_n1466), .B2 (CLOCK_slo__sro_n1468));
INV_X1 CLOCK_slo__xsl_c1060 (.ZN (CLOCK_slo__xsl_n1441), .A (n_11));
AND2_X2 CLOCK_slo__xsl_c1063 (.ZN (n_11), .A1 (slo__sro_n247), .A2 (slo__sro_n248));
XNOR2_X1 CLOCK_slo__sro_c1105 (.ZN (p_1[3]), .A (CLOCK_slo__sro_n1465), .B (n_3));
INV_X1 slo__sro_c602 (.ZN (slo__sro_n834), .A (n_18));
NAND2_X1 slo__sro_c603 (.ZN (slo__sro_n833), .A1 (p_0[18]), .A2 (Multiplier[18]));
NOR2_X1 slo__sro_c604 (.ZN (slo__sro_n832), .A1 (p_0[18]), .A2 (Multiplier[18]));
OAI21_X1 slo__sro_c605 (.ZN (n_19), .A (slo__sro_n833), .B1 (slo__sro_n834), .B2 (slo__sro_n832));
XNOR2_X1 slo__sro_c606 (.ZN (slo__sro_n831), .A (p_0[18]), .B (Multiplier[18]));
XNOR2_X1 slo__sro_c607 (.ZN (p_1[18]), .A (slo__sro_n831), .B (n_18));
NOR2_X1 CLOCK_slo__sro_c1129 (.ZN (CLOCK_slo__sro_n1494), .A1 (n_5), .A2 (Multiplier[5]));
OAI21_X1 CLOCK_slo__sro_c1130 (.ZN (n_6), .A (CLOCK_slo__sro_n1495), .B1 (CLOCK_slo__sro_n1496), .B2 (CLOCK_slo__sro_n1494));
XNOR2_X1 CLOCK_slo__sro_c1131 (.ZN (CLOCK_slo__sro_n1493), .A (n_5), .B (Multiplier[5]));
XNOR2_X1 CLOCK_slo__sro_c1132 (.ZN (p_1[5]), .A (CLOCK_slo__sro_n1493), .B (p_0[5]));
OR2_X1 CLOCK_slo__sro_c1283 (.ZN (CLOCK_slo__sro_n1660), .A1 (p_0[30]), .A2 (n_34));
INV_X1 CLOCK_slo__xsl_c1196 (.ZN (CLOCK_slo__xsl_n1562), .A (n_9));
INV_X1 CLOCK_slo__xsl_c1197 (.ZN (CLOCK_slo__xsl_n1561), .A (CLOCK_slo__xsl_n1562));
OAI22_X1 CLOCK_slo__sro_c1284 (.ZN (n_31), .A1 (n_32), .A2 (CLOCK_slo__sro_n1660)
    , .B1 (CLOCK_slo__sro_n1661), .B2 (n_30));
NAND2_X1 CLOCK_slo__sro_c1241 (.ZN (CLOCK_slo__sro_n1616), .A1 (p_0[12]), .A2 (Multiplier[12]));
OAI21_X1 CLOCK_slo__sro_c1242 (.ZN (CLOCK_slo__sro_n1615), .A (slo__sro_n133), .B1 (p_0[12]), .B2 (Multiplier[12]));
NAND2_X1 CLOCK_slo__sro_c1243 (.ZN (CLOCK_slo__sro_n1614), .A1 (CLOCK_slo__sro_n1615), .A2 (CLOCK_slo__sro_n1616));
XNOR2_X1 CLOCK_slo__sro_c1244 (.ZN (CLOCK_slo__sro_n1613), .A (p_0[12]), .B (Multiplier[12]));
XNOR2_X1 CLOCK_slo__sro_c1245 (.ZN (p_1[12]), .A (CLOCK_slo__sro_n1613), .B (slo__sro_n133));

endmodule //datapath__0_171

module datapath__0_167 (p_0, p_1, p_2);

output [31:0] p_2;
input [31:0] p_0;
input [31:0] p_1;
wire slo__sro_n759;
wire CLOCK_slo__sro_n1331;
wire slo__sro_n703;
wire n_1;
wire n_2;
wire n_3;
wire n_4;
wire n_6;
wire slo__sro_n996;
wire n_10;
wire n_11;
wire n_12;
wire n_13;
wire n_14;
wire n_16;
wire n_17;
wire n_18;
wire n_19;
wire n_21;
wire n_22;
wire n_23;
wire n_24;
wire n_25;
wire n_26;
wire n_27;
wire n_28;
wire n_29;
wire n_30;
wire n_32;
wire n_0;
wire n_34;
wire n_33;
wire CLOCK_slo__sro_n1335;
wire slo__sro_n67;
wire slo__sro_n68;
wire slo__sro_n69;
wire slo__sro_n70;
wire slo__sro_n156;
wire slo__sro_n157;
wire slo__sro_n158;
wire slo__sro_n159;
wire slo__sro_n104;
wire slo__sro_n105;
wire slo__sro_n106;
wire slo__sro_n107;
wire slo__sro_n171;
wire slo__sro_n172;
wire slo__sro_n173;
wire slo__sro_n174;
wire slo__sro_n184;
wire slo__sro_n185;
wire slo__sro_n186;
wire slo__sro_n187;
wire slo__sro_n188;
wire slo__sro_n205;
wire slo__sro_n206;
wire slo__sro_n228;
wire slo__sro_n229;
wire slo__sro_n230;
wire slo__sro_n231;
wire slo__sro_n232;
wire slo__sro_n275;
wire slo__sro_n276;
wire slo__sro_n277;
wire slo__sro_n278;
wire slo__sro_n337;
wire slo__sro_n338;
wire slo__sro_n339;
wire slo__sro_n340;
wire slo__sro_n341;
wire slo__sro_n342;
wire slo__sro_n467;
wire slo__sro_n468;
wire slo__sro_n469;
wire slo__sro_n470;
wire slo__sro_n471;
wire slo__sro_n487;
wire slo__sro_n488;
wire slo__sro_n489;
wire slo__sro_n490;
wire slo__sro_n704;
wire slo__sro_n705;
wire slo__sro_n706;
wire CLOCK_slo__mro_n1726;
wire slo__sro_n544;
wire slo__sro_n545;
wire slo__sro_n546;
wire slo__sro_n547;
wire slo__sro_n760;
wire slo__sro_n761;
wire slo__sro_n762;
wire slo__sro_n798;
wire slo__sro_n799;
wire slo__sro_n800;
wire slo__sro_n801;
wire slo__sro_n802;
wire slo__sro_n997;
wire slo__sro_n998;
wire slo__sro_n999;
wire slo__sro_n1000;
wire CLOCK_slo__sro_n1332;
wire CLOCK_slo__sro_n1333;
wire CLOCK_slo__sro_n1334;
wire CLOCK_slo__sro_n1369;
wire CLOCK_slo__sro_n1370;
wire CLOCK_slo__sro_n1371;
wire CLOCK_slo__mro_n1703;


INV_X1 i_36 (.ZN (n_34), .A (p_0[30]));
INV_X1 i_35 (.ZN (n_33), .A (p_1[30]));
INV_X2 i_34 (.ZN (n_32), .A (n_30));
XNOR2_X1 CLOCK_slo__mro_c876 (.ZN (p_2[16]), .A (n_16), .B (slo__sro_n544));
XOR2_X1 i_32 (.Z (p_2[31]), .A (p_0[31]), .B (slo__sro_n996));
OAI22_X1 i_31 (.ZN (n_0), .A1 (n_34), .A2 (p_1[30]), .B1 (p_0[30]), .B2 (n_33));
XNOR2_X1 i_0 (.ZN (p_2[30]), .A (n_32), .B (n_0));
FA_X1 i_30 (.CO (n_30), .S (p_2[29]), .A (p_0[29]), .B (p_1[29]), .CI (n_29));
FA_X1 i_29 (.CO (n_29), .S (p_2[28]), .A (p_0[28]), .B (p_1[28]), .CI (n_28));
FA_X1 i_28 (.CO (n_28), .S (p_2[27]), .A (p_0[27]), .B (p_1[27]), .CI (n_27));
INV_X1 slo__sro_c168 (.ZN (slo__sro_n232), .A (n_19));
INV_X1 slo__sro_c98 (.ZN (slo__sro_n159), .A (n_23));
FA_X1 i_25 (.CO (n_25), .S (p_2[24]), .A (p_0[24]), .B (p_1[24]), .CI (n_24));
INV_X1 slo__sro_c112 (.ZN (slo__sro_n174), .A (n_3));
FA_X1 i_23 (.CO (n_23), .S (p_2[22]), .A (p_0[22]), .B (p_1[22]), .CI (n_22));
FA_X1 i_22 (.CO (n_22), .S (p_2[21]), .A (p_0[21]), .B (p_1[21]), .CI (n_21));
FA_X1 i_21 (.CO (n_21), .S (p_2[20]), .A (p_0[20]), .B (p_1[20]), .CI (slo__sro_n229));
INV_X1 slo__sro_c210 (.ZN (slo__sro_n278), .A (p_1[9]));
NAND2_X1 slo__sro_c357 (.ZN (slo__sro_n470), .A1 (n_4), .A2 (p_0[4]));
FA_X1 i_18 (.CO (n_18), .S (p_2[17]), .A (p_0[17]), .B (p_1[17]), .CI (n_17));
NAND2_X1 slo__sro_c533 (.ZN (slo__sro_n761), .A1 (p_1[2]), .A2 (p_0[2]));
FA_X1 i_16 (.CO (n_16), .S (p_2[15]), .A (p_0[15]), .B (p_1[15]), .CI (CLOCK_slo__sro_n1332));
NAND2_X1 CLOCK_slo__sro_c950 (.ZN (CLOCK_slo__sro_n1371), .A1 (n_10), .A2 (p_0[10]));
FA_X1 i_14 (.CO (n_14), .S (p_2[13]), .A (p_0[13]), .B (p_1[13]), .CI (n_13));
NAND2_X1 slo__sro_c113 (.ZN (slo__sro_n173), .A1 (p_1[3]), .A2 (p_0[3]));
FA_X1 i_12 (.CO (n_12), .S (p_2[11]), .A (p_0[11]), .B (p_1[11]), .CI (n_11));
INV_X1 slo__sro_c486 (.ZN (slo__sro_n706), .A (p_1[5]));
NAND2_X1 slo__sro_c143 (.ZN (slo__sro_n206), .A1 (n_26), .A2 (p_0[26]));
INV_X1 slo__sro_c698 (.ZN (slo__sro_n1000), .A (n_30));
NAND2_X1 slo__sro_c487 (.ZN (slo__sro_n705), .A1 (slo__sro_n468), .A2 (p_0[5]));
INV_X1 slo__sro_c532 (.ZN (slo__sro_n762), .A (n_2));
INV_X1 slo__sro_c372 (.ZN (slo__sro_n490), .A (n_6));
INV_X1 slo__sro_c126 (.ZN (slo__sro_n188), .A (slo__sro_n799));
INV_X1 slo__sro_c561 (.ZN (slo__sro_n802), .A (p_1[7]));
FA_X1 i_2 (.CO (n_2), .S (p_2[1]), .A (p_0[1]), .B (p_1[1]), .CI (n_1));
HA_X1 i_1 (.CO (n_1), .S (p_2[0]), .A (p_0[0]), .B (p_1[0]));
INV_X2 slo__sro_c5 (.ZN (slo__sro_n70), .A (n_25));
NAND2_X1 slo__sro_c6 (.ZN (slo__sro_n69), .A1 (p_1[25]), .A2 (p_0[25]));
NOR2_X1 slo__sro_c7 (.ZN (slo__sro_n68), .A1 (p_1[25]), .A2 (p_0[25]));
OAI21_X2 slo__sro_c8 (.ZN (n_26), .A (slo__sro_n69), .B1 (slo__sro_n70), .B2 (slo__sro_n68));
XNOR2_X1 slo__sro_c9 (.ZN (slo__sro_n67), .A (p_1[25]), .B (p_0[25]));
XNOR2_X1 slo__sro_c10 (.ZN (p_2[25]), .A (slo__sro_n67), .B (n_25));
NAND2_X1 slo__sro_c99 (.ZN (slo__sro_n158), .A1 (p_1[23]), .A2 (p_0[23]));
NOR2_X1 slo__sro_c100 (.ZN (slo__sro_n157), .A1 (p_1[23]), .A2 (p_0[23]));
OAI21_X1 slo__sro_c101 (.ZN (n_24), .A (slo__sro_n158), .B1 (slo__sro_n159), .B2 (slo__sro_n157));
XNOR2_X1 slo__sro_c102 (.ZN (slo__sro_n156), .A (p_1[23]), .B (p_0[23]));
XNOR2_X1 slo__sro_c103 (.ZN (p_2[23]), .A (slo__sro_n156), .B (n_23));
INV_X1 slo__sro_c45 (.ZN (slo__sro_n107), .A (n_12));
NAND2_X1 slo__sro_c46 (.ZN (slo__sro_n106), .A1 (p_1[12]), .A2 (p_0[12]));
NOR2_X1 slo__sro_c47 (.ZN (slo__sro_n105), .A1 (p_1[12]), .A2 (p_0[12]));
OAI21_X1 slo__sro_c48 (.ZN (n_13), .A (slo__sro_n106), .B1 (slo__sro_n107), .B2 (slo__sro_n105));
XNOR2_X1 slo__sro_c49 (.ZN (slo__sro_n104), .A (p_1[12]), .B (p_0[12]));
XNOR2_X1 slo__sro_c50 (.ZN (p_2[12]), .A (slo__sro_n104), .B (n_12));
NOR2_X1 slo__sro_c114 (.ZN (slo__sro_n172), .A1 (p_1[3]), .A2 (p_0[3]));
OAI21_X1 slo__sro_c115 (.ZN (n_4), .A (slo__sro_n173), .B1 (slo__sro_n174), .B2 (slo__sro_n172));
XNOR2_X2 slo__sro_c116 (.ZN (slo__sro_n171), .A (p_1[3]), .B (p_0[3]));
XNOR2_X2 slo__sro_c117 (.ZN (p_2[3]), .A (slo__sro_n171), .B (n_3));
NAND2_X1 slo__sro_c127 (.ZN (slo__sro_n187), .A1 (p_1[8]), .A2 (p_0[8]));
NOR2_X1 slo__sro_c128 (.ZN (slo__sro_n186), .A1 (p_1[8]), .A2 (p_0[8]));
OAI21_X2 slo__sro_c129 (.ZN (slo__sro_n185), .A (slo__sro_n187), .B1 (slo__sro_n186), .B2 (slo__sro_n188));
XNOR2_X1 slo__sro_c130 (.ZN (slo__sro_n184), .A (p_1[8]), .B (p_0[8]));
XNOR2_X1 slo__sro_c131 (.ZN (p_2[8]), .A (slo__sro_n184), .B (slo__sro_n799));
OAI21_X1 slo__sro_c144 (.ZN (slo__sro_n205), .A (p_1[26]), .B1 (n_26), .B2 (p_0[26]));
NAND2_X1 slo__sro_c145 (.ZN (n_27), .A1 (slo__sro_n205), .A2 (slo__sro_n206));
INV_X1 CLOCK_slo__sro_c917 (.ZN (CLOCK_slo__sro_n1335), .A (n_14));
NAND2_X1 CLOCK_slo__sro_c918 (.ZN (CLOCK_slo__sro_n1334), .A1 (p_1[14]), .A2 (p_0[14]));
NAND2_X1 slo__sro_c169 (.ZN (slo__sro_n231), .A1 (p_1[19]), .A2 (p_0[19]));
NOR2_X1 slo__sro_c170 (.ZN (slo__sro_n230), .A1 (p_1[19]), .A2 (p_0[19]));
OAI21_X1 slo__sro_c171 (.ZN (slo__sro_n229), .A (slo__sro_n231), .B1 (slo__sro_n232), .B2 (slo__sro_n230));
XNOR2_X1 slo__sro_c172 (.ZN (slo__sro_n228), .A (p_1[19]), .B (p_0[19]));
XNOR2_X1 slo__sro_c173 (.ZN (p_2[19]), .A (slo__sro_n228), .B (n_19));
NAND2_X1 slo__sro_c211 (.ZN (slo__sro_n277), .A1 (slo__sro_n185), .A2 (p_0[9]));
NOR2_X2 slo__sro_c212 (.ZN (slo__sro_n276), .A1 (slo__sro_n185), .A2 (p_0[9]));
OAI21_X2 slo__sro_c213 (.ZN (n_10), .A (slo__sro_n277), .B1 (slo__sro_n276), .B2 (slo__sro_n278));
XNOR2_X1 slo__sro_c214 (.ZN (slo__sro_n275), .A (slo__sro_n185), .B (p_0[9]));
XNOR2_X1 slo__sro_c215 (.ZN (p_2[9]), .A (slo__sro_n275), .B (p_1[9]));
INV_X1 slo__sro_c356 (.ZN (slo__sro_n471), .A (p_1[4]));
INV_X1 slo__sro_c242 (.ZN (slo__sro_n342), .A (p_0[18]));
INV_X1 slo__sro_c243 (.ZN (slo__sro_n341), .A (p_1[18]));
NAND2_X1 slo__sro_c244 (.ZN (slo__sro_n340), .A1 (p_1[18]), .A2 (p_0[18]));
NAND2_X1 slo__sro_c245 (.ZN (slo__sro_n339), .A1 (slo__sro_n341), .A2 (slo__sro_n342));
NAND2_X1 slo__sro_c246 (.ZN (slo__sro_n338), .A1 (n_18), .A2 (slo__sro_n339));
NAND2_X2 slo__sro_c247 (.ZN (n_19), .A1 (slo__sro_n338), .A2 (slo__sro_n340));
XNOR2_X1 slo__sro_c248 (.ZN (slo__sro_n337), .A (p_1[18]), .B (p_0[18]));
XNOR2_X1 slo__sro_c249 (.ZN (p_2[18]), .A (n_18), .B (slo__sro_n337));
NOR2_X1 slo__sro_c358 (.ZN (slo__sro_n469), .A1 (n_4), .A2 (p_0[4]));
OAI21_X1 slo__sro_c359 (.ZN (slo__sro_n468), .A (slo__sro_n470), .B1 (slo__sro_n471), .B2 (slo__sro_n469));
XNOR2_X1 slo__sro_c360 (.ZN (slo__sro_n467), .A (n_4), .B (p_0[4]));
XNOR2_X1 slo__sro_c361 (.ZN (p_2[4]), .A (p_1[4]), .B (slo__sro_n467));
NAND2_X1 slo__sro_c373 (.ZN (slo__sro_n489), .A1 (p_1[6]), .A2 (p_0[6]));
NOR2_X2 slo__sro_c374 (.ZN (slo__sro_n488), .A1 (p_1[6]), .A2 (p_0[6]));
NOR2_X1 slo__sro_c488 (.ZN (slo__sro_n704), .A1 (slo__sro_n468), .A2 (p_0[5]));
OAI21_X1 slo__sro_c489 (.ZN (n_6), .A (slo__sro_n705), .B1 (slo__sro_n706), .B2 (slo__sro_n704));
XNOR2_X1 slo__sro_c490 (.ZN (slo__sro_n703), .A (slo__sro_n468), .B (p_0[5]));
XNOR2_X1 slo__sro_c491 (.ZN (p_2[5]), .A (slo__sro_n703), .B (p_1[5]));
INV_X1 slo__sro_c422 (.ZN (slo__sro_n547), .A (n_16));
NAND2_X1 slo__sro_c423 (.ZN (slo__sro_n546), .A1 (p_1[16]), .A2 (p_0[16]));
NOR2_X1 slo__sro_c424 (.ZN (slo__sro_n545), .A1 (p_1[16]), .A2 (p_0[16]));
OAI21_X1 slo__sro_c425 (.ZN (n_17), .A (slo__sro_n546), .B1 (slo__sro_n547), .B2 (slo__sro_n545));
XNOR2_X1 slo__sro_c426 (.ZN (slo__sro_n544), .A (p_1[16]), .B (p_0[16]));
XNOR2_X1 CLOCK_slo__mro_c1292 (.ZN (CLOCK_slo__mro_n1726), .A (n_6), .B (p_0[6]));
NOR2_X1 slo__sro_c534 (.ZN (slo__sro_n760), .A1 (p_1[2]), .A2 (p_0[2]));
OAI21_X2 slo__sro_c535 (.ZN (n_3), .A (slo__sro_n761), .B1 (slo__sro_n762), .B2 (slo__sro_n760));
XNOR2_X2 slo__sro_c536 (.ZN (slo__sro_n759), .A (p_1[2]), .B (p_0[2]));
XNOR2_X2 slo__sro_c537 (.ZN (p_2[2]), .A (slo__sro_n759), .B (n_2));
NAND2_X1 slo__sro_c562 (.ZN (slo__sro_n801), .A1 (slo__sro_n487), .A2 (p_0[7]));
NOR2_X1 slo__sro_c563 (.ZN (slo__sro_n800), .A1 (slo__sro_n487), .A2 (p_0[7]));
OAI21_X2 slo__sro_c564 (.ZN (slo__sro_n799), .A (slo__sro_n801), .B1 (slo__sro_n802), .B2 (slo__sro_n800));
XNOR2_X2 slo__sro_c565 (.ZN (slo__sro_n798), .A (slo__sro_n487), .B (p_0[7]));
XNOR2_X2 slo__sro_c566 (.ZN (p_2[7]), .A (slo__sro_n798), .B (p_1[7]));
NOR2_X1 slo__sro_c699 (.ZN (slo__sro_n999), .A1 (n_33), .A2 (p_0[30]));
NAND2_X1 slo__sro_c700 (.ZN (slo__sro_n998), .A1 (slo__sro_n999), .A2 (slo__sro_n1000));
OR2_X1 slo__sro_c701 (.ZN (slo__sro_n997), .A1 (p_1[30]), .A2 (n_34));
OAI21_X1 slo__sro_c702 (.ZN (slo__sro_n996), .A (slo__sro_n998), .B1 (n_32), .B2 (slo__sro_n997));
XNOR2_X1 CLOCK_slo__mro_c1293 (.ZN (p_2[6]), .A (CLOCK_slo__mro_n1726), .B (p_1[6]));
NOR2_X1 CLOCK_slo__sro_c919 (.ZN (CLOCK_slo__sro_n1333), .A1 (p_1[14]), .A2 (p_0[14]));
OAI21_X1 CLOCK_slo__sro_c920 (.ZN (CLOCK_slo__sro_n1332), .A (CLOCK_slo__sro_n1334)
    , .B1 (CLOCK_slo__sro_n1335), .B2 (CLOCK_slo__sro_n1333));
XNOR2_X1 CLOCK_slo__sro_c921 (.ZN (CLOCK_slo__sro_n1331), .A (p_1[14]), .B (p_0[14]));
XNOR2_X1 CLOCK_slo__sro_c922 (.ZN (p_2[14]), .A (CLOCK_slo__sro_n1331), .B (n_14));
OAI21_X2 CLOCK_slo__sro_c951 (.ZN (CLOCK_slo__sro_n1370), .A (p_1[10]), .B1 (n_10), .B2 (p_0[10]));
NAND2_X1 CLOCK_slo__sro_c952 (.ZN (n_11), .A1 (CLOCK_slo__sro_n1370), .A2 (CLOCK_slo__sro_n1371));
XNOR2_X1 CLOCK_slo__sro_c953 (.ZN (CLOCK_slo__sro_n1369), .A (n_10), .B (p_0[10]));
XNOR2_X1 CLOCK_slo__sro_c954 (.ZN (p_2[10]), .A (CLOCK_slo__sro_n1369), .B (p_1[10]));
OAI21_X2 CLOCK_slo__sro_c972 (.ZN (slo__sro_n487), .A (slo__sro_n489), .B1 (slo__sro_n488), .B2 (slo__sro_n490));
XNOR2_X1 CLOCK_slo__mro_c1259 (.ZN (p_2[26]), .A (CLOCK_slo__mro_n1703), .B (n_26));
XNOR2_X1 CLOCK_slo__mro_c1258 (.ZN (CLOCK_slo__mro_n1703), .A (p_1[26]), .B (p_0[26]));

endmodule //datapath__0_167

module datapath__0_166 (drc_ipoPP_0, Multiplier, p_0, p_1);

output [31:0] p_1;
input [31:0] Multiplier;
input [31:0] p_0;
input drc_ipoPP_0;
wire CLOCK_slo__sro_n1757;
wire n_1;
wire n_2;
wire n_3;
wire n_4;
wire n_5;
wire n_6;
wire n_8;
wire n_9;
wire n_10;
wire n_12;
wire n_15;
wire n_16;
wire n_17;
wire n_18;
wire n_19;
wire n_20;
wire n_21;
wire n_22;
wire n_23;
wire n_24;
wire n_25;
wire n_26;
wire n_28;
wire n_29;
wire n_30;
wire n_32;
wire n_0;
wire n_34;
wire n_33;
wire slo__sro_n59;
wire slo__sro_n60;
wire slo__sro_n61;
wire slo__sro_n62;
wire slo__sro_n72;
wire slo__sro_n73;
wire slo__sro_n74;
wire slo__sro_n75;
wire slo__sro_n85;
wire slo__sro_n86;
wire slo__sro_n87;
wire slo__sro_n88;
wire slo__sro_n89;
wire slo__sro_n119;
wire slo__sro_n120;
wire slo__sro_n121;
wire slo__sro_n122;
wire slo__sro_n134;
wire slo__sro_n135;
wire slo__sro_n136;
wire slo__sro_n137;
wire slo__sro_n138;
wire slo__sro_n151;
wire slo__sro_n152;
wire slo__sro_n153;
wire slo__sro_n154;
wire slo__sro_n166;
wire slo__sro_n167;
wire slo__sro_n168;
wire slo__sro_n185;
wire slo__sro_n186;
wire slo__sro_n187;
wire slo__sro_n188;
wire CLOCK_slo__sro_n1758;
wire slo__sro_n212;
wire slo__sro_n213;
wire slo__sro_n214;
wire slo__sro_n230;
wire slo__sro_n231;
wire slo__sro_n232;
wire slo__sro_n233;
wire slo__sro_n440;
wire slo__sro_n441;
wire slo__sro_n442;
wire slo__sro_n443;
wire slo__sro_n741;
wire slo__sro_n742;
wire slo__sro_n743;
wire slo__sro_n744;
wire slo__sro_n745;
wire slo__sro_n808;
wire slo__sro_n809;
wire slo__sro_n810;
wire slo__sro_n811;
wire CLOCK_slo__sro_n1117;
wire CLOCK_slo__sro_n1118;
wire CLOCK_slo__sro_n1119;
wire CLOCK_slo__sro_n1120;
wire CLOCK_slo__mro_n1679;
wire CLOCK_slo__sro_n1229;
wire CLOCK_slo__sro_n1230;
wire CLOCK_slo__sro_n1231;
wire CLOCK_slo__sro_n1232;
wire CLOCK_slo__sro_n1233;
wire CLOCK_slo__sro_n1314;
wire CLOCK_slo__sro_n1315;
wire CLOCK_slo__sro_n1316;
wire CLOCK_slo__sro_n1317;
wire CLOCK_slo__sro_n1756;
wire CLOCK_slo__sro_n1561;
wire CLOCK_slo__sro_n1562;
wire CLOCK_slo__sro_n1563;
wire CLOCK_slo__sro_n1759;
wire CLOCK_slo__sro_n1799;
wire CLOCK_slo__sro_n1800;
wire CLOCK_slo__sro_n1801;
wire CLOCK_slo__sro_n1802;
wire CLOCK_slo__sro_n1803;


INV_X1 i_36 (.ZN (n_34), .A (Multiplier[30]));
INV_X1 i_35 (.ZN (n_33), .A (p_0[30]));
INV_X1 i_34 (.ZN (n_32), .A (n_30));
XOR2_X1 i_32 (.Z (p_1[31]), .A (Multiplier[31]), .B (CLOCK_slo__sro_n1799));
OAI22_X1 i_31 (.ZN (n_0), .A1 (n_34), .A2 (p_0[30]), .B1 (Multiplier[30]), .B2 (n_33));
XNOR2_X1 i_0 (.ZN (p_1[30]), .A (n_32), .B (n_0));
FA_X1 i_30 (.CO (n_30), .S (p_1[29]), .A (Multiplier[29]), .B (p_0[29]), .CI (n_29));
FA_X1 i_29 (.CO (n_29), .S (p_1[28]), .A (Multiplier[28]), .B (p_0[28]), .CI (n_28));
INV_X1 slo__sro_c126 (.ZN (slo__sro_n188), .A (n_20));
INV_X2 slo__sro_c61 (.ZN (slo__sro_n122), .A (slo__sro_n135));
INV_X1 slo__sro_c29 (.ZN (slo__sro_n89), .A (p_0[26]));
FA_X1 i_25 (.CO (n_25), .S (p_1[24]), .A (Multiplier[24]), .B (p_0[24]), .CI (n_24));
NAND2_X1 slo__sro_c105 (.ZN (slo__sro_n168), .A1 (Multiplier[27]), .A2 (slo__sro_n86));
FA_X1 i_23 (.CO (n_23), .S (p_1[22]), .A (Multiplier[22]), .B (p_0[22]), .CI (n_22));
NOR2_X2 CLOCK_slo__sro_c1464 (.ZN (CLOCK_slo__sro_n1757), .A1 (p_0[7]), .A2 (Multiplier[7]));
NAND2_X1 slo__sro_c153 (.ZN (slo__sro_n214), .A1 (Multiplier[12]), .A2 (p_0[12]));
FA_X1 i_20 (.CO (n_20), .S (p_1[19]), .A (Multiplier[19]), .B (p_0[19]), .CI (n_19));
FA_X1 i_19 (.CO (n_19), .S (p_1[18]), .A (Multiplier[18]), .B (p_0[18]), .CI (n_18));
INV_X2 slo__sro_c15 (.ZN (slo__sro_n75), .A (n_25));
NOR2_X1 slo__sro_c575 (.ZN (slo__sro_n743), .A1 (p_0[13]), .A2 (Multiplier[13]));
FA_X1 i_16 (.CO (n_16), .S (p_1[15]), .A (Multiplier[15]), .B (p_0[15]), .CI (n_15));
INV_X1 CLOCK_slo__sro_c1462 (.ZN (CLOCK_slo__sro_n1759), .A (CLOCK_slo__sro_n1230));
INV_X1 slo__sro_c632 (.ZN (slo__sro_n811), .A (n_2));
INV_X1 slo__sro_c169 (.ZN (slo__sro_n233), .A (n_9));
INV_X1 slo__sro_c77 (.ZN (slo__sro_n138), .A (n_10));
INV_X1 slo__sro_c91 (.ZN (slo__sro_n154), .A (n_23));
INV_X1 slo__sro_c573 (.ZN (slo__sro_n745), .A (slo__sro_n212));
FA_X1 i_9 (.CO (n_9), .S (p_1[8]), .A (Multiplier[8]), .B (p_0[8]), .CI (n_8));
INV_X1 CLOCK_slo__sro_c1504 (.ZN (CLOCK_slo__sro_n1803), .A (n_30));
INV_X1 CLOCK_slo__sro_c1031 (.ZN (CLOCK_slo__sro_n1317), .A (slo__sro_n742));
FA_X1 i_6 (.CO (n_6), .S (p_1[5]), .A (Multiplier[5]), .B (p_0[5]), .CI (n_5));
XNOR2_X2 CLOCK_slo__mro_c1381 (.ZN (p_1[12]), .A (CLOCK_slo__mro_n1679), .B (n_12));
FA_X1 i_4 (.CO (n_4), .S (p_1[3]), .A (Multiplier[3]), .B (p_0[3]), .CI (n_3));
INV_X1 CLOCK_slo__sro_c839 (.ZN (CLOCK_slo__sro_n1120), .A (p_0[4]));
FA_X1 i_2 (.CO (n_2), .S (p_1[1]), .A (Multiplier[1]), .B (p_0[1]), .CI (n_1));
HA_X1 i_1 (.CO (n_1), .S (p_1[0]), .A (Multiplier[0]), .B (p_0[0]));
INV_X1 slo__sro_c1 (.ZN (slo__sro_n62), .A (n_17));
NAND2_X1 slo__sro_c2 (.ZN (slo__sro_n61), .A1 (p_0[17]), .A2 (Multiplier[17]));
NOR2_X1 slo__sro_c3 (.ZN (slo__sro_n60), .A1 (p_0[17]), .A2 (Multiplier[17]));
OAI21_X1 slo__sro_c4 (.ZN (n_18), .A (slo__sro_n61), .B1 (slo__sro_n62), .B2 (slo__sro_n60));
XNOR2_X1 slo__sro_c5 (.ZN (slo__sro_n59), .A (p_0[17]), .B (Multiplier[17]));
XNOR2_X1 slo__sro_c6 (.ZN (p_1[17]), .A (slo__sro_n59), .B (n_17));
NAND2_X1 slo__sro_c16 (.ZN (slo__sro_n74), .A1 (p_0[25]), .A2 (Multiplier[25]));
NOR2_X1 slo__sro_c17 (.ZN (slo__sro_n73), .A1 (p_0[25]), .A2 (Multiplier[25]));
OAI21_X2 slo__sro_c18 (.ZN (n_26), .A (slo__sro_n74), .B1 (slo__sro_n75), .B2 (slo__sro_n73));
XNOR2_X2 slo__sro_c19 (.ZN (slo__sro_n72), .A (p_0[25]), .B (Multiplier[25]));
XNOR2_X2 slo__sro_c20 (.ZN (p_1[25]), .A (slo__sro_n72), .B (n_25));
NAND2_X1 slo__sro_c30 (.ZN (slo__sro_n88), .A1 (n_26), .A2 (Multiplier[26]));
NOR2_X1 slo__sro_c31 (.ZN (slo__sro_n87), .A1 (n_26), .A2 (Multiplier[26]));
OAI21_X2 slo__sro_c32 (.ZN (slo__sro_n86), .A (slo__sro_n88), .B1 (slo__sro_n89), .B2 (slo__sro_n87));
XNOR2_X2 slo__sro_c33 (.ZN (slo__sro_n85), .A (n_26), .B (Multiplier[26]));
XNOR2_X2 slo__sro_c34 (.ZN (p_1[26]), .A (slo__sro_n85), .B (p_0[26]));
NAND2_X1 slo__sro_c62 (.ZN (slo__sro_n121), .A1 (p_0[11]), .A2 (Multiplier[11]));
NOR2_X1 slo__sro_c63 (.ZN (slo__sro_n120), .A1 (p_0[11]), .A2 (Multiplier[11]));
OAI21_X2 slo__sro_c64 (.ZN (n_12), .A (slo__sro_n121), .B1 (slo__sro_n120), .B2 (slo__sro_n122));
XNOR2_X1 slo__sro_c65 (.ZN (slo__sro_n119), .A (p_0[11]), .B (drc_ipoPP_0));
XNOR2_X1 slo__sro_c66 (.ZN (p_1[11]), .A (slo__sro_n119), .B (slo__sro_n135));
NAND2_X1 slo__sro_c78 (.ZN (slo__sro_n137), .A1 (p_0[10]), .A2 (Multiplier[10]));
NOR2_X1 slo__sro_c79 (.ZN (slo__sro_n136), .A1 (p_0[10]), .A2 (Multiplier[10]));
OAI21_X2 slo__sro_c80 (.ZN (slo__sro_n135), .A (slo__sro_n137), .B1 (slo__sro_n136), .B2 (slo__sro_n138));
XNOR2_X1 slo__sro_c81 (.ZN (slo__sro_n134), .A (p_0[10]), .B (Multiplier[10]));
XNOR2_X2 slo__sro_c82 (.ZN (p_1[10]), .A (n_10), .B (slo__sro_n134));
NAND2_X1 slo__sro_c92 (.ZN (slo__sro_n153), .A1 (p_0[23]), .A2 (Multiplier[23]));
NOR2_X1 slo__sro_c93 (.ZN (slo__sro_n152), .A1 (p_0[23]), .A2 (Multiplier[23]));
OAI21_X1 slo__sro_c94 (.ZN (n_24), .A (slo__sro_n153), .B1 (slo__sro_n154), .B2 (slo__sro_n152));
XNOR2_X1 slo__sro_c95 (.ZN (slo__sro_n151), .A (p_0[23]), .B (Multiplier[23]));
XNOR2_X1 slo__sro_c96 (.ZN (p_1[23]), .A (slo__sro_n151), .B (n_23));
OAI21_X1 slo__sro_c106 (.ZN (slo__sro_n167), .A (p_0[27]), .B1 (slo__sro_n86), .B2 (Multiplier[27]));
NAND2_X1 slo__sro_c107 (.ZN (n_28), .A1 (slo__sro_n167), .A2 (slo__sro_n168));
XNOR2_X2 slo__sro_c108 (.ZN (slo__sro_n166), .A (slo__sro_n86), .B (Multiplier[27]));
XNOR2_X2 slo__sro_c109 (.ZN (p_1[27]), .A (slo__sro_n166), .B (p_0[27]));
NAND2_X1 slo__sro_c127 (.ZN (slo__sro_n187), .A1 (p_0[20]), .A2 (Multiplier[20]));
NOR2_X1 slo__sro_c128 (.ZN (slo__sro_n186), .A1 (p_0[20]), .A2 (Multiplier[20]));
OAI21_X1 slo__sro_c129 (.ZN (n_21), .A (slo__sro_n187), .B1 (slo__sro_n188), .B2 (slo__sro_n186));
XNOR2_X1 slo__sro_c130 (.ZN (slo__sro_n185), .A (p_0[20]), .B (Multiplier[20]));
XNOR2_X1 slo__sro_c131 (.ZN (p_1[20]), .A (slo__sro_n185), .B (n_20));
OAI21_X1 slo__sro_c154 (.ZN (slo__sro_n213), .A (n_12), .B1 (p_0[12]), .B2 (Multiplier[12]));
NAND2_X1 slo__sro_c155 (.ZN (slo__sro_n212), .A1 (slo__sro_n213), .A2 (slo__sro_n214));
OAI21_X1 CLOCK_slo__sro_c1243 (.ZN (CLOCK_slo__sro_n1562), .A (n_21), .B1 (p_0[21]), .B2 (Multiplier[21]));
XNOR2_X1 CLOCK_slo__sro_c1466 (.ZN (CLOCK_slo__sro_n1756), .A (p_0[7]), .B (Multiplier[7]));
NAND2_X1 slo__sro_c170 (.ZN (slo__sro_n232), .A1 (p_0[9]), .A2 (Multiplier[9]));
NOR2_X1 slo__sro_c171 (.ZN (slo__sro_n231), .A1 (p_0[9]), .A2 (Multiplier[9]));
OAI21_X2 slo__sro_c172 (.ZN (n_10), .A (slo__sro_n232), .B1 (slo__sro_n233), .B2 (slo__sro_n231));
XNOR2_X1 slo__sro_c173 (.ZN (slo__sro_n230), .A (p_0[9]), .B (Multiplier[9]));
XNOR2_X1 slo__sro_c174 (.ZN (p_1[9]), .A (slo__sro_n230), .B (n_9));
NAND2_X1 slo__sro_c574 (.ZN (slo__sro_n744), .A1 (p_0[13]), .A2 (Multiplier[13]));
INV_X1 slo__sro_c325 (.ZN (slo__sro_n443), .A (n_16));
NAND2_X1 slo__sro_c326 (.ZN (slo__sro_n442), .A1 (p_0[16]), .A2 (Multiplier[16]));
NOR2_X1 slo__sro_c327 (.ZN (slo__sro_n441), .A1 (p_0[16]), .A2 (Multiplier[16]));
OAI21_X1 slo__sro_c328 (.ZN (n_17), .A (slo__sro_n442), .B1 (slo__sro_n443), .B2 (slo__sro_n441));
XNOR2_X1 slo__sro_c329 (.ZN (slo__sro_n440), .A (p_0[16]), .B (Multiplier[16]));
XNOR2_X1 slo__sro_c330 (.ZN (p_1[16]), .A (slo__sro_n440), .B (n_16));
OAI21_X2 slo__sro_c576 (.ZN (slo__sro_n742), .A (slo__sro_n744), .B1 (slo__sro_n743), .B2 (slo__sro_n745));
XNOR2_X1 slo__sro_c577 (.ZN (slo__sro_n741), .A (p_0[13]), .B (Multiplier[13]));
XNOR2_X1 slo__sro_c578 (.ZN (p_1[13]), .A (slo__sro_n741), .B (slo__sro_n212));
NAND2_X1 slo__sro_c633 (.ZN (slo__sro_n810), .A1 (p_0[2]), .A2 (Multiplier[2]));
NOR2_X1 slo__sro_c634 (.ZN (slo__sro_n809), .A1 (p_0[2]), .A2 (Multiplier[2]));
OAI21_X1 slo__sro_c635 (.ZN (n_3), .A (slo__sro_n810), .B1 (slo__sro_n809), .B2 (slo__sro_n811));
XNOR2_X1 slo__sro_c636 (.ZN (slo__sro_n808), .A (p_0[2]), .B (Multiplier[2]));
XNOR2_X1 slo__sro_c637 (.ZN (p_1[2]), .A (slo__sro_n808), .B (n_2));
NAND2_X1 CLOCK_slo__sro_c840 (.ZN (CLOCK_slo__sro_n1119), .A1 (n_4), .A2 (Multiplier[4]));
NOR2_X1 CLOCK_slo__sro_c841 (.ZN (CLOCK_slo__sro_n1118), .A1 (n_4), .A2 (Multiplier[4]));
OAI21_X1 CLOCK_slo__sro_c842 (.ZN (n_5), .A (CLOCK_slo__sro_n1119), .B1 (CLOCK_slo__sro_n1120), .B2 (CLOCK_slo__sro_n1118));
XNOR2_X1 CLOCK_slo__sro_c843 (.ZN (CLOCK_slo__sro_n1117), .A (n_4), .B (Multiplier[4]));
XNOR2_X1 CLOCK_slo__sro_c844 (.ZN (p_1[4]), .A (CLOCK_slo__sro_n1117), .B (p_0[4]));
XNOR2_X2 CLOCK_slo__mro_c1380 (.ZN (CLOCK_slo__mro_n1679), .A (p_0[12]), .B (Multiplier[12]));
INV_X1 CLOCK_slo__sro_c954 (.ZN (CLOCK_slo__sro_n1233), .A (n_6));
NAND2_X1 CLOCK_slo__sro_c955 (.ZN (CLOCK_slo__sro_n1232), .A1 (p_0[6]), .A2 (Multiplier[6]));
NOR2_X1 CLOCK_slo__sro_c956 (.ZN (CLOCK_slo__sro_n1231), .A1 (p_0[6]), .A2 (Multiplier[6]));
OAI21_X1 CLOCK_slo__sro_c957 (.ZN (CLOCK_slo__sro_n1230), .A (CLOCK_slo__sro_n1232)
    , .B1 (CLOCK_slo__sro_n1231), .B2 (CLOCK_slo__sro_n1233));
XNOR2_X1 CLOCK_slo__sro_c958 (.ZN (CLOCK_slo__sro_n1229), .A (p_0[6]), .B (Multiplier[6]));
XNOR2_X1 CLOCK_slo__sro_c959 (.ZN (p_1[6]), .A (CLOCK_slo__sro_n1229), .B (n_6));
NAND2_X1 CLOCK_slo__sro_c1032 (.ZN (CLOCK_slo__sro_n1316), .A1 (p_0[14]), .A2 (Multiplier[14]));
NOR2_X1 CLOCK_slo__sro_c1033 (.ZN (CLOCK_slo__sro_n1315), .A1 (p_0[14]), .A2 (Multiplier[14]));
OAI21_X1 CLOCK_slo__sro_c1034 (.ZN (n_15), .A (CLOCK_slo__sro_n1316), .B1 (CLOCK_slo__sro_n1317), .B2 (CLOCK_slo__sro_n1315));
XNOR2_X1 CLOCK_slo__sro_c1035 (.ZN (CLOCK_slo__sro_n1314), .A (p_0[14]), .B (Multiplier[14]));
XNOR2_X1 CLOCK_slo__sro_c1036 (.ZN (p_1[14]), .A (CLOCK_slo__sro_n1314), .B (slo__sro_n742));
NAND2_X1 CLOCK_slo__sro_c1463 (.ZN (CLOCK_slo__sro_n1758), .A1 (p_0[7]), .A2 (Multiplier[7]));
NAND2_X1 CLOCK_slo__sro_c1242 (.ZN (CLOCK_slo__sro_n1563), .A1 (p_0[21]), .A2 (Multiplier[21]));
NAND2_X1 CLOCK_slo__sro_c1244 (.ZN (n_22), .A1 (CLOCK_slo__sro_n1563), .A2 (CLOCK_slo__sro_n1562));
XNOR2_X2 CLOCK_slo__sro_c1245 (.ZN (CLOCK_slo__sro_n1561), .A (p_0[21]), .B (Multiplier[21]));
XNOR2_X2 CLOCK_slo__sro_c1246 (.ZN (p_1[21]), .A (CLOCK_slo__sro_n1561), .B (n_21));
OAI21_X2 CLOCK_slo__sro_c1465 (.ZN (n_8), .A (CLOCK_slo__sro_n1758), .B1 (CLOCK_slo__sro_n1759), .B2 (CLOCK_slo__sro_n1757));
XNOR2_X1 CLOCK_slo__sro_c1467 (.ZN (p_1[7]), .A (CLOCK_slo__sro_n1756), .B (CLOCK_slo__sro_n1230));
NOR2_X1 CLOCK_slo__sro_c1505 (.ZN (CLOCK_slo__sro_n1802), .A1 (n_33), .A2 (Multiplier[30]));
NAND2_X1 CLOCK_slo__sro_c1506 (.ZN (CLOCK_slo__sro_n1801), .A1 (CLOCK_slo__sro_n1802), .A2 (CLOCK_slo__sro_n1803));
OR2_X1 CLOCK_slo__sro_c1507 (.ZN (CLOCK_slo__sro_n1800), .A1 (p_0[30]), .A2 (n_34));
OAI21_X1 CLOCK_slo__sro_c1508 (.ZN (CLOCK_slo__sro_n1799), .A (CLOCK_slo__sro_n1801)
    , .B1 (n_32), .B2 (CLOCK_slo__sro_n1800));

endmodule //datapath__0_166

module datapath__0_162 (drc_ipoPP_0, p_0_19_PP_0, p_0, p_1, p_2);

output [31:0] p_2;
input [31:0] p_0;
input [31:0] p_1;
input drc_ipoPP_0;
input p_0_19_PP_0;
wire n_1;
wire n_2;
wire n_4;
wire n_6;
wire n_7;
wire n_8;
wire n_9;
wire n_10;
wire n_11;
wire n_12;
wire n_14;
wire n_16;
wire n_17;
wire n_18;
wire n_19;
wire n_20;
wire n_21;
wire n_22;
wire n_23;
wire n_24;
wire n_26;
wire n_28;
wire n_29;
wire n_30;
wire n_32;
wire n_0;
wire n_34;
wire n_33;
wire n_31;
wire slo__sro_n76;
wire slo__sro_n77;
wire slo__sro_n78;
wire slo__sro_n79;
wire slo__sro_n104;
wire slo__sro_n105;
wire slo__sro_n106;
wire slo__sro_n107;
wire slo__sro_n119;
wire slo__sro_n120;
wire slo__sro_n121;
wire slo__sro_n122;
wire slo__sro_n123;
wire slo__sro_n148;
wire slo__sro_n149;
wire slo__sro_n150;
wire slo__sro_n151;
wire slo__sro_n163;
wire slo__sro_n164;
wire slo__sro_n165;
wire slo__sro_n166;
wire slo__sro_n167;
wire slo__sro_n446;
wire slo__sro_n447;
wire slo__sro_n448;
wire slo__sro_n222;
wire slo__sro_n223;
wire slo__sro_n224;
wire slo__sro_n225;
wire slo__sro_n610;
wire slo__sro_n611;
wire slo__sro_n612;
wire slo__sro_n613;
wire slo__mro_n623;
wire slo__sro_n641;
wire slo__sro_n642;
wire slo__sro_n643;
wire slo__sro_n644;
wire slo__sro_n669;
wire slo__sro_n670;
wire slo__sro_n671;
wire slo__sro_n672;
wire slo__sro_n673;
wire slo__sro_n688;
wire slo__sro_n689;
wire slo__sro_n690;
wire slo__sro_n705;
wire slo__sro_n706;
wire slo__sro_n707;
wire slo__sro_n708;
wire slo__n838;
wire CLOCK_slo__sro_n1012;
wire CLOCK_slo__sro_n1013;
wire CLOCK_slo__sro_n1014;
wire CLOCK_slo__sro_n1015;
wire CLOCK_slo__sro_n1016;
wire CLOCK_slo__sro_n1040;
wire CLOCK_slo__sro_n1041;
wire CLOCK_slo__sro_n1042;
wire CLOCK_slo__sro_n1043;
wire CLOCK_slo__sro_n1044;
wire CLOCK_slo__sro_n1075;
wire CLOCK_slo__sro_n1076;
wire CLOCK_slo__sro_n1077;
wire CLOCK_slo__sro_n1078;
wire CLOCK_slo__sro_n1079;
wire CLOCK_slo__sro_n1080;
wire CLOCK_slo__sro_n1221;
wire CLOCK_slo__sro_n1222;
wire CLOCK_slo__sro_n1223;
wire CLOCK_slo__sro_n1224;
wire CLOCK_slo__sro_n1240;
wire CLOCK_slo__sro_n1241;
wire CLOCK_slo__sro_n1242;
wire CLOCK_slo__sro_n1243;
wire CLOCK_slo__sro_n1244;
wire CLOCK_slo__sro_n1245;


INV_X1 i_36 (.ZN (n_34), .A (p_0[30]));
INV_X1 i_35 (.ZN (n_33), .A (p_1[30]));
INV_X1 i_34 (.ZN (n_32), .A (n_30));
OAI33_X1 i_33 (.ZN (n_31), .A1 (n_34), .A2 (p_1[30]), .A3 (n_32), .B1 (p_0[30]), .B2 (n_33), .B3 (n_30));
XOR2_X1 i_32 (.Z (p_2[31]), .A (p_0[31]), .B (n_31));
OAI22_X1 i_31 (.ZN (n_0), .A1 (n_34), .A2 (p_1[30]), .B1 (p_0[30]), .B2 (n_33));
XNOR2_X1 i_0 (.ZN (p_2[30]), .A (n_32), .B (n_0));
INV_X1 slo__sro_c57 (.ZN (slo__sro_n123), .A (n_24));
FA_X1 i_29 (.CO (n_29), .S (p_2[28]), .A (p_0[28]), .B (p_1[28]), .CI (n_28));
FA_X1 i_28 (.CO (n_28), .S (p_2[27]), .A (p_0[27]), .B (p_1[27]), .CI (CLOCK_slo__sro_n1013));
FA_X1 i_26 (.CO (n_26), .S (p_2[25]), .A (p_0[25]), .B (p_1[25]), .CI (slo__sro_n120));
INV_X1 slo__sro_c84 (.ZN (slo__sro_n151), .A (n_19));
XNOR2_X2 slo__mro_c478 (.ZN (slo__mro_n623), .A (p_1[2]), .B (p_0[2]));
INV_X1 slo__sro_c43 (.ZN (slo__sro_n107), .A (n_29));
INV_X1 CLOCK_slo__sro_c921 (.ZN (CLOCK_slo__sro_n1245), .A (p_0[11]));
FA_X1 i_21 (.CO (n_21), .S (p_2[20]), .A (p_0[20]), .B (p_1[20]), .CI (n_20));
INV_X1 slo__sro_c98 (.ZN (slo__sro_n167), .A (n_14));
FA_X1 i_17 (.CO (n_17), .S (p_2[16]), .A (p_0[16]), .B (p_1[16]), .CI (n_16));
FA_X1 i_16 (.CO (n_16), .S (p_2[15]), .A (p_0[15]), .B (p_1[15]), .CI (slo__sro_n164));
INV_X1 slo__sro_c459 (.ZN (slo__sro_n613), .A (n_23));
FA_X1 i_14 (.CO (n_14), .S (p_2[13]), .A (p_0[13]), .B (p_1[13]), .CI (CLOCK_slo__sro_n1041));
INV_X1 CLOCK_slo__sro_c792 (.ZN (CLOCK_slo__sro_n1080), .A (p_0[17]));
XNOR2_X1 slo__sro_c336 (.ZN (p_2[2]), .A (slo__mro_n623), .B (n_2));
INV_X1 slo__sro_c514 (.ZN (slo__sro_n673), .A (p_1[4]));
FA_X1 i_9 (.CO (n_9), .S (p_2[8]), .A (p_0[8]), .B (p_1[8]), .CI (n_8));
FA_X1 i_8 (.CO (n_8), .S (p_2[7]), .A (p_0[7]), .B (p_1[7]), .CI (n_7));
FA_X1 i_7 (.CO (n_7), .S (p_2[6]), .A (p_0[6]), .B (p_1[6]), .CI (n_6));
FA_X1 i_6 (.CO (n_6), .S (p_2[5]), .A (p_0[5]), .B (p_1[5]), .CI (slo__sro_n670));
INV_X1 slo__sro_c544 (.ZN (slo__sro_n708), .A (n_18));
NAND2_X1 slo__sro_c460 (.ZN (slo__sro_n612), .A1 (p_1[23]), .A2 (p_0[23]));
FA_X1 i_2 (.CO (n_2), .S (p_2[1]), .A (p_0[1]), .B (p_1[1]), .CI (n_1));
HA_X1 i_1 (.CO (n_1), .S (p_2[0]), .A (p_0[0]), .B (p_1[0]));
INV_X1 slo__sro_c14 (.ZN (slo__sro_n79), .A (n_22));
NAND2_X1 slo__sro_c15 (.ZN (slo__sro_n78), .A1 (p_1[22]), .A2 (p_0[22]));
NOR2_X1 slo__sro_c16 (.ZN (slo__sro_n77), .A1 (p_1[22]), .A2 (p_0[22]));
OAI21_X2 slo__sro_c17 (.ZN (n_23), .A (slo__sro_n78), .B1 (slo__sro_n79), .B2 (slo__sro_n77));
XNOR2_X1 slo__sro_c18 (.ZN (slo__sro_n76), .A (p_1[22]), .B (drc_ipoPP_0));
XNOR2_X1 slo__sro_c19 (.ZN (p_2[22]), .A (slo__sro_n76), .B (n_22));
NAND2_X1 slo__sro_c44 (.ZN (slo__sro_n106), .A1 (p_1[29]), .A2 (p_0[29]));
NOR2_X1 slo__sro_c45 (.ZN (slo__sro_n105), .A1 (p_1[29]), .A2 (p_0[29]));
OAI21_X1 slo__sro_c46 (.ZN (n_30), .A (slo__sro_n106), .B1 (slo__sro_n107), .B2 (slo__sro_n105));
XNOR2_X1 slo__sro_c47 (.ZN (slo__sro_n104), .A (p_1[29]), .B (p_0[29]));
XNOR2_X1 slo__sro_c48 (.ZN (p_2[29]), .A (n_29), .B (slo__sro_n104));
NAND2_X1 slo__sro_c58 (.ZN (slo__sro_n122), .A1 (p_1[24]), .A2 (p_0[24]));
NOR2_X2 slo__sro_c59 (.ZN (slo__sro_n121), .A1 (p_1[24]), .A2 (p_0[24]));
OAI21_X1 slo__sro_c60 (.ZN (slo__sro_n120), .A (slo__sro_n122), .B1 (slo__sro_n123), .B2 (slo__sro_n121));
XNOR2_X1 slo__sro_c61 (.ZN (slo__sro_n119), .A (p_1[24]), .B (p_0[24]));
XNOR2_X1 slo__sro_c62 (.ZN (p_2[24]), .A (slo__sro_n119), .B (n_24));
NAND2_X1 slo__sro_c85 (.ZN (slo__sro_n150), .A1 (p_1[19]), .A2 (p_0[19]));
NOR2_X1 slo__sro_c86 (.ZN (slo__sro_n149), .A1 (p_1[19]), .A2 (p_0[19]));
OAI21_X1 slo__sro_c87 (.ZN (n_20), .A (slo__sro_n150), .B1 (slo__sro_n151), .B2 (slo__sro_n149));
XNOR2_X1 slo__sro_c88 (.ZN (slo__sro_n148), .A (p_1[19]), .B (p_0_19_PP_0));
XNOR2_X1 slo__sro_c89 (.ZN (p_2[19]), .A (n_19), .B (slo__sro_n148));
NAND2_X1 slo__sro_c99 (.ZN (slo__sro_n166), .A1 (p_1[14]), .A2 (p_0[14]));
NOR2_X1 slo__sro_c100 (.ZN (slo__sro_n165), .A1 (p_1[14]), .A2 (p_0[14]));
OAI21_X1 slo__sro_c101 (.ZN (slo__sro_n164), .A (slo__sro_n166), .B1 (slo__sro_n167), .B2 (slo__sro_n165));
XNOR2_X1 slo__sro_c102 (.ZN (slo__sro_n163), .A (p_1[14]), .B (p_0[14]));
XNOR2_X1 slo__sro_c103 (.ZN (p_2[14]), .A (slo__sro_n163), .B (n_14));
NAND2_X1 slo__sro_c332 (.ZN (slo__sro_n448), .A1 (p_1[2]), .A2 (p_0[2]));
NOR2_X2 slo__sro_c333 (.ZN (slo__sro_n447), .A1 (p_1[2]), .A2 (p_0[2]));
OAI21_X2 slo__sro_c334 (.ZN (slo__sro_n446), .A (slo__sro_n448), .B1 (slo__sro_n447), .B2 (slo__n838));
INV_X1 slo__sro_c151 (.ZN (slo__sro_n225), .A (n_10));
NAND2_X1 slo__sro_c152 (.ZN (slo__sro_n224), .A1 (p_1[10]), .A2 (p_0[10]));
NOR2_X1 slo__sro_c153 (.ZN (slo__sro_n223), .A1 (p_1[10]), .A2 (p_0[10]));
OAI21_X1 slo__sro_c154 (.ZN (n_11), .A (slo__sro_n224), .B1 (slo__sro_n225), .B2 (slo__sro_n223));
XNOR2_X1 slo__sro_c155 (.ZN (slo__sro_n222), .A (p_1[10]), .B (p_0[10]));
XNOR2_X1 slo__sro_c156 (.ZN (p_2[10]), .A (slo__sro_n222), .B (n_10));
NOR2_X1 slo__sro_c461 (.ZN (slo__sro_n611), .A1 (p_1[23]), .A2 (p_0[23]));
OAI21_X2 slo__sro_c462 (.ZN (n_24), .A (slo__sro_n612), .B1 (slo__sro_n611), .B2 (slo__sro_n613));
XNOR2_X1 slo__sro_c463 (.ZN (slo__sro_n610), .A (p_1[23]), .B (p_0[23]));
XNOR2_X2 slo__sro_c464 (.ZN (p_2[23]), .A (slo__sro_n610), .B (n_23));
INV_X1 slo__sro_c494 (.ZN (slo__sro_n644), .A (n_9));
NAND2_X1 slo__sro_c495 (.ZN (slo__sro_n643), .A1 (p_1[9]), .A2 (p_0[9]));
NOR2_X1 slo__sro_c496 (.ZN (slo__sro_n642), .A1 (p_1[9]), .A2 (p_0[9]));
OAI21_X1 slo__sro_c497 (.ZN (n_10), .A (slo__sro_n643), .B1 (slo__sro_n644), .B2 (slo__sro_n642));
XNOR2_X1 slo__sro_c498 (.ZN (slo__sro_n641), .A (p_1[9]), .B (p_0[9]));
XNOR2_X2 slo__sro_c499 (.ZN (p_2[9]), .A (n_9), .B (slo__sro_n641));
NAND2_X1 slo__sro_c515 (.ZN (slo__sro_n672), .A1 (n_4), .A2 (p_0[4]));
NOR2_X1 slo__sro_c516 (.ZN (slo__sro_n671), .A1 (n_4), .A2 (p_0[4]));
OAI21_X1 slo__sro_c517 (.ZN (slo__sro_n670), .A (slo__sro_n672), .B1 (slo__sro_n671), .B2 (slo__sro_n673));
XNOR2_X1 slo__sro_c518 (.ZN (slo__sro_n669), .A (n_4), .B (p_0[4]));
XNOR2_X1 slo__sro_c519 (.ZN (p_2[4]), .A (slo__sro_n669), .B (p_1[4]));
NAND2_X1 slo__sro_c529 (.ZN (slo__sro_n690), .A1 (slo__sro_n446), .A2 (p_0[3]));
OAI21_X1 slo__sro_c530 (.ZN (slo__sro_n689), .A (p_1[3]), .B1 (slo__sro_n446), .B2 (p_0[3]));
NAND2_X2 slo__sro_c531 (.ZN (n_4), .A1 (slo__sro_n689), .A2 (slo__sro_n690));
XNOR2_X2 slo__sro_c532 (.ZN (slo__sro_n688), .A (slo__sro_n446), .B (p_0[3]));
XNOR2_X1 slo__sro_c533 (.ZN (p_2[3]), .A (slo__sro_n688), .B (p_1[3]));
NAND2_X1 slo__sro_c545 (.ZN (slo__sro_n707), .A1 (p_1[18]), .A2 (p_0[18]));
NOR2_X1 slo__sro_c546 (.ZN (slo__sro_n706), .A1 (p_1[18]), .A2 (p_0[18]));
OAI21_X1 slo__sro_c547 (.ZN (n_19), .A (slo__sro_n707), .B1 (slo__sro_n708), .B2 (slo__sro_n706));
XNOR2_X1 slo__sro_c548 (.ZN (slo__sro_n705), .A (p_1[18]), .B (p_0[18]));
XNOR2_X1 slo__sro_c549 (.ZN (p_2[18]), .A (n_18), .B (slo__sro_n705));
INV_X1 slo__L1_c633 (.ZN (slo__n838), .A (n_2));
INV_X1 CLOCK_slo__sro_c731 (.ZN (CLOCK_slo__sro_n1016), .A (n_26));
NAND2_X1 CLOCK_slo__sro_c732 (.ZN (CLOCK_slo__sro_n1015), .A1 (p_1[26]), .A2 (p_0[26]));
NOR2_X1 CLOCK_slo__sro_c733 (.ZN (CLOCK_slo__sro_n1014), .A1 (p_1[26]), .A2 (p_0[26]));
OAI21_X1 CLOCK_slo__sro_c734 (.ZN (CLOCK_slo__sro_n1013), .A (CLOCK_slo__sro_n1015)
    , .B1 (CLOCK_slo__sro_n1014), .B2 (CLOCK_slo__sro_n1016));
XNOR2_X1 CLOCK_slo__sro_c735 (.ZN (CLOCK_slo__sro_n1012), .A (p_1[26]), .B (p_0[26]));
XNOR2_X1 CLOCK_slo__sro_c736 (.ZN (p_2[26]), .A (CLOCK_slo__sro_n1012), .B (n_26));
INV_X1 CLOCK_slo__sro_c756 (.ZN (CLOCK_slo__sro_n1044), .A (n_12));
NAND2_X1 CLOCK_slo__sro_c757 (.ZN (CLOCK_slo__sro_n1043), .A1 (p_1[12]), .A2 (p_0[12]));
NOR2_X1 CLOCK_slo__sro_c758 (.ZN (CLOCK_slo__sro_n1042), .A1 (p_1[12]), .A2 (p_0[12]));
OAI21_X1 CLOCK_slo__sro_c759 (.ZN (CLOCK_slo__sro_n1041), .A (CLOCK_slo__sro_n1043)
    , .B1 (CLOCK_slo__sro_n1044), .B2 (CLOCK_slo__sro_n1042));
XNOR2_X1 CLOCK_slo__sro_c760 (.ZN (CLOCK_slo__sro_n1040), .A (p_1[12]), .B (p_0[12]));
XNOR2_X1 CLOCK_slo__sro_c761 (.ZN (p_2[12]), .A (CLOCK_slo__sro_n1040), .B (n_12));
INV_X1 CLOCK_slo__sro_c793 (.ZN (CLOCK_slo__sro_n1079), .A (p_1[17]));
NAND2_X1 CLOCK_slo__sro_c794 (.ZN (CLOCK_slo__sro_n1078), .A1 (p_1[17]), .A2 (p_0[17]));
NAND2_X1 CLOCK_slo__sro_c795 (.ZN (CLOCK_slo__sro_n1077), .A1 (CLOCK_slo__sro_n1079), .A2 (CLOCK_slo__sro_n1080));
NAND2_X1 CLOCK_slo__sro_c796 (.ZN (CLOCK_slo__sro_n1076), .A1 (n_17), .A2 (CLOCK_slo__sro_n1077));
NAND2_X1 CLOCK_slo__sro_c797 (.ZN (n_18), .A1 (CLOCK_slo__sro_n1076), .A2 (CLOCK_slo__sro_n1078));
XNOR2_X1 CLOCK_slo__sro_c798 (.ZN (CLOCK_slo__sro_n1075), .A (p_1[17]), .B (p_0[17]));
XNOR2_X1 CLOCK_slo__sro_c799 (.ZN (p_2[17]), .A (n_17), .B (CLOCK_slo__sro_n1075));
INV_X1 CLOCK_slo__sro_c903 (.ZN (CLOCK_slo__sro_n1224), .A (n_21));
NAND2_X1 CLOCK_slo__sro_c904 (.ZN (CLOCK_slo__sro_n1223), .A1 (p_1[21]), .A2 (p_0[21]));
NOR2_X1 CLOCK_slo__sro_c905 (.ZN (CLOCK_slo__sro_n1222), .A1 (p_1[21]), .A2 (p_0[21]));
OAI21_X2 CLOCK_slo__sro_c906 (.ZN (n_22), .A (CLOCK_slo__sro_n1223), .B1 (CLOCK_slo__sro_n1224), .B2 (CLOCK_slo__sro_n1222));
XNOR2_X1 CLOCK_slo__sro_c907 (.ZN (CLOCK_slo__sro_n1221), .A (p_1[21]), .B (p_0[21]));
XNOR2_X1 CLOCK_slo__sro_c908 (.ZN (p_2[21]), .A (CLOCK_slo__sro_n1221), .B (n_21));
INV_X1 CLOCK_slo__sro_c922 (.ZN (CLOCK_slo__sro_n1244), .A (p_1[11]));
NAND2_X1 CLOCK_slo__sro_c923 (.ZN (CLOCK_slo__sro_n1243), .A1 (p_1[11]), .A2 (p_0[11]));
NAND2_X1 CLOCK_slo__sro_c924 (.ZN (CLOCK_slo__sro_n1242), .A1 (CLOCK_slo__sro_n1244), .A2 (CLOCK_slo__sro_n1245));
NAND2_X1 CLOCK_slo__sro_c925 (.ZN (CLOCK_slo__sro_n1241), .A1 (n_11), .A2 (CLOCK_slo__sro_n1242));
NAND2_X1 CLOCK_slo__sro_c926 (.ZN (n_12), .A1 (CLOCK_slo__sro_n1241), .A2 (CLOCK_slo__sro_n1243));
XNOR2_X1 CLOCK_slo__sro_c927 (.ZN (CLOCK_slo__sro_n1240), .A (p_1[11]), .B (p_0[11]));
XNOR2_X1 CLOCK_slo__sro_c928 (.ZN (p_2[11]), .A (n_11), .B (CLOCK_slo__sro_n1240));

endmodule //datapath__0_162

module datapath__0_161 (drc_ipoPP_0, Multiplier, p_0, p_1);

output [31:0] p_1;
input [31:0] Multiplier;
input [31:0] p_0;
input drc_ipoPP_0;
wire CLOCK_slo__sro_n1600;
wire CLOCK_slo__sro_n1598;
wire n_1;
wire n_2;
wire n_3;
wire n_4;
wire n_6;
wire n_7;
wire n_8;
wire n_9;
wire n_10;
wire n_12;
wire n_13;
wire n_14;
wire n_15;
wire n_16;
wire n_17;
wire n_18;
wire n_19;
wire n_20;
wire n_21;
wire n_22;
wire n_23;
wire n_26;
wire n_27;
wire n_28;
wire n_30;
wire n_32;
wire n_0;
wire n_34;
wire n_33;
wire n_31;
wire slo__sro_n59;
wire slo__sro_n60;
wire slo__sro_n61;
wire slo__sro_n62;
wire CLOCK_slo__sro_n1100;
wire slo__sro_n73;
wire slo__sro_n74;
wire slo__sro_n75;
wire slo__sro_n76;
wire slo__sro_n89;
wire slo__sro_n90;
wire slo__sro_n91;
wire slo__sro_n92;
wire slo__n843;
wire slo__sro_n105;
wire slo__sro_n106;
wire slo__sro_n107;
wire slo__sro_n133;
wire slo__sro_n134;
wire slo__sro_n135;
wire slo__sro_n136;
wire slo__sro_n168;
wire slo__sro_n169;
wire slo__sro_n170;
wire slo__sro_n171;
wire slo__sro_n213;
wire slo__sro_n214;
wire slo__sro_n215;
wire slo__sro_n216;
wire slo__sro_n255;
wire slo__sro_n256;
wire slo__sro_n257;
wire slo__sro_n268;
wire slo__sro_n269;
wire slo__sro_n270;
wire slo__sro_n271;
wire slo__sro_n272;
wire slo__sro_n445;
wire slo__sro_n446;
wire slo__sro_n447;
wire CLOCK_slo__sro_n1597;
wire slo__sro_n658;
wire slo__sro_n659;
wire slo__sro_n660;
wire slo__sro_n661;
wire slo__sro_n765;
wire slo__sro_n766;
wire slo__sro_n767;
wire slo__sro_n768;
wire slo__mro_n786;
wire slo__sro_n825;
wire slo__sro_n826;
wire slo__sro_n827;
wire slo__sro_n828;
wire CLOCK_slo__sro_n1064;
wire CLOCK_slo__sro_n1065;
wire CLOCK_slo__sro_n1066;
wire CLOCK_slo__sro_n1067;
wire CLOCK_slo__sro_n1068;
wire CLOCK_slo__mro_n1081;
wire CLOCK_slo__sro_n1101;
wire CLOCK_slo__sro_n1102;
wire CLOCK_slo__sro_n1103;
wire CLOCK_slo__mro_n1162;
wire CLOCK_slo__sro_n1206;
wire CLOCK_slo__sro_n1207;
wire CLOCK_slo__sro_n1208;
wire CLOCK_slo__sro_n1209;
wire CLOCK_slo__sro_n1210;
wire CLOCK_slo__sro_n1233;
wire CLOCK_slo__sro_n1234;
wire CLOCK_slo__sro_n1235;
wire CLOCK_slo__sro_n1236;
wire CLOCK_slo__sro_n1599;
wire CLOCK_slo__sro_n1449;
wire CLOCK_slo__sro_n1450;
wire CLOCK_slo__sro_n1451;
wire CLOCK_slo__sro_n1452;


INV_X1 i_36 (.ZN (n_34), .A (Multiplier[30]));
INV_X1 i_35 (.ZN (n_33), .A (p_0[30]));
INV_X1 i_34 (.ZN (n_32), .A (n_30));
OAI33_X1 i_33 (.ZN (n_31), .A1 (n_34), .A2 (p_0[30]), .A3 (n_32), .B1 (Multiplier[30])
    , .B2 (n_33), .B3 (n_30));
XOR2_X1 i_32 (.Z (p_1[31]), .A (Multiplier[31]), .B (n_31));
OAI22_X1 i_31 (.ZN (n_0), .A1 (n_34), .A2 (p_0[30]), .B1 (Multiplier[30]), .B2 (n_33));
XNOR2_X1 i_0 (.ZN (p_1[30]), .A (n_32), .B (n_0));
INV_X1 slo__sro_c145 (.ZN (slo__sro_n216), .A (p_0[14]));
INV_X1 slo__sro_c103 (.ZN (slo__sro_n171), .A (slo__sro_n133));
XNOR2_X1 CLOCK_slo__sro_c1389 (.ZN (CLOCK_slo__sro_n1597), .A (p_0[11]), .B (Multiplier[11]));
FA_X1 i_27 (.CO (n_27), .S (p_1[26]), .A (Multiplier[26]), .B (p_0[26]), .CI (n_26));
FA_X1 i_26 (.CO (n_26), .S (p_1[25]), .A (Multiplier[25]), .B (p_0[25]), .CI (slo__sro_n73));
INV_X1 slo__sro_c29 (.ZN (slo__sro_n92), .A (n_20));
XNOR2_X2 CLOCK_slo__mro_c857 (.ZN (CLOCK_slo__mro_n1081), .A (CLOCK_slo__sro_n1065), .B (Multiplier[24]));
FA_X1 i_23 (.CO (n_23), .S (p_1[22]), .A (Multiplier[22]), .B (p_0[22]), .CI (n_22));
INV_X1 slo__sro_c589 (.ZN (slo__sro_n768), .A (n_12));
INV_X1 slo__sro_c45 (.ZN (slo__sro_n107), .A (n_19));
INV_X1 slo__sro_c72 (.ZN (slo__sro_n136), .A (n_28));
INV_X1 CLOCK_slo__sro_c1385 (.ZN (CLOCK_slo__sro_n1600), .A (slo__sro_n269));
INV_X1 slo__sro_c525 (.ZN (slo__sro_n661), .A (p_0[21]));
XNOR2_X2 CLOCK_slo__mro_c937 (.ZN (CLOCK_slo__mro_n1162), .A (p_0[28]), .B (Multiplier[28]));
INV_X1 slo__sro_c197 (.ZN (slo__sro_n272), .A (n_10));
NAND2_X1 slo__sro_c185 (.ZN (slo__sro_n257), .A1 (n_15), .A2 (Multiplier[15]));
INV_X1 slo__sro_c15 (.ZN (slo__sro_n76), .A (CLOCK_slo__sro_n1065));
XNOR2_X2 slo__mro_c609 (.ZN (slo__mro_n786), .A (n_19), .B (drc_ipoPP_0));
NAND2_X1 CLOCK_slo__sro_c1386 (.ZN (CLOCK_slo__sro_n1599), .A1 (p_0[11]), .A2 (Multiplier[11]));
FA_X1 i_10 (.CO (n_10), .S (p_1[9]), .A (Multiplier[9]), .B (p_0[9]), .CI (n_9));
OAI21_X1 CLOCK_slo__sro_c1388 (.ZN (n_12), .A (CLOCK_slo__sro_n1599), .B1 (CLOCK_slo__sro_n1600), .B2 (CLOCK_slo__sro_n1598));
FA_X1 i_8 (.CO (n_8), .S (p_1[7]), .A (Multiplier[7]), .B (p_0[7]), .CI (n_7));
FA_X1 i_7 (.CO (n_7), .S (p_1[6]), .A (Multiplier[6]), .B (p_0[6]), .CI (n_6));
FA_X1 i_6 (.CO (n_6), .S (p_1[5]), .A (Multiplier[5]), .B (p_0[5]), .CI (CLOCK_slo__sro_n1207));
INV_X1 CLOCK_slo__sro_c1015 (.ZN (CLOCK_slo__sro_n1236), .A (n_8));
FA_X1 i_4 (.CO (n_4), .S (p_1[3]), .A (Multiplier[3]), .B (p_0[3]), .CI (n_3));
FA_X1 i_3 (.CO (n_3), .S (p_1[2]), .A (Multiplier[2]), .B (p_0[2]), .CI (n_2));
FA_X1 i_2 (.CO (n_2), .S (p_1[1]), .A (Multiplier[1]), .B (p_0[1]), .CI (n_1));
HA_X1 i_1 (.CO (n_1), .S (p_1[0]), .A (Multiplier[0]), .B (p_0[0]));
INV_X1 slo__sro_c1 (.ZN (slo__sro_n62), .A (n_13));
NAND2_X1 slo__sro_c2 (.ZN (slo__sro_n61), .A1 (p_0[13]), .A2 (Multiplier[13]));
NOR2_X2 slo__sro_c3 (.ZN (slo__sro_n60), .A1 (p_0[13]), .A2 (Multiplier[13]));
OAI21_X1 CLOCK_slo__sro_c1230 (.ZN (n_28), .A (CLOCK_slo__sro_n1451), .B1 (CLOCK_slo__sro_n1452), .B2 (CLOCK_slo__sro_n1450));
XNOR2_X1 slo__sro_c5 (.ZN (slo__sro_n59), .A (p_0[13]), .B (Multiplier[13]));
XNOR2_X1 slo__sro_c6 (.ZN (p_1[13]), .A (slo__sro_n59), .B (n_13));
NAND2_X1 slo__sro_c16 (.ZN (slo__sro_n75), .A1 (p_0[24]), .A2 (Multiplier[24]));
NOR2_X2 slo__sro_c17 (.ZN (slo__sro_n74), .A1 (p_0[24]), .A2 (Multiplier[24]));
OAI21_X1 slo__sro_c18 (.ZN (slo__sro_n73), .A (slo__sro_n75), .B1 (slo__sro_n74), .B2 (slo__sro_n76));
INV_X1 CLOCK_slo__sro_c876 (.ZN (CLOCK_slo__sro_n1103), .A (n_16));
NAND2_X1 CLOCK_slo__sro_c877 (.ZN (CLOCK_slo__sro_n1102), .A1 (p_0[16]), .A2 (Multiplier[16]));
NAND2_X1 slo__sro_c30 (.ZN (slo__sro_n91), .A1 (p_0[20]), .A2 (Multiplier[20]));
NOR2_X1 slo__sro_c31 (.ZN (slo__sro_n90), .A1 (p_0[20]), .A2 (Multiplier[20]));
OAI21_X1 slo__sro_c32 (.ZN (n_21), .A (slo__sro_n91), .B1 (slo__sro_n90), .B2 (slo__sro_n92));
XNOR2_X1 slo__sro_c33 (.ZN (slo__sro_n89), .A (p_0[20]), .B (Multiplier[20]));
XNOR2_X1 slo__sro_c34 (.ZN (p_1[20]), .A (slo__sro_n89), .B (n_20));
NAND2_X1 slo__sro_c46 (.ZN (slo__sro_n106), .A1 (p_0[19]), .A2 (Multiplier[19]));
NOR2_X1 slo__sro_c47 (.ZN (slo__sro_n105), .A1 (p_0[19]), .A2 (Multiplier[19]));
OAI21_X1 slo__sro_c48 (.ZN (n_20), .A (slo__sro_n106), .B1 (slo__sro_n107), .B2 (slo__sro_n105));
INV_X1 slo__L1_c661 (.ZN (slo__n843), .A (n_17));
NAND2_X1 CLOCK_slo__sro_c844 (.ZN (CLOCK_slo__sro_n1067), .A1 (p_0[23]), .A2 (Multiplier[23]));
NAND2_X1 slo__sro_c73 (.ZN (slo__sro_n135), .A1 (p_0[28]), .A2 (Multiplier[28]));
NOR2_X1 slo__sro_c74 (.ZN (slo__sro_n134), .A1 (p_0[28]), .A2 (Multiplier[28]));
OAI21_X1 slo__sro_c75 (.ZN (slo__sro_n133), .A (slo__sro_n135), .B1 (slo__sro_n136), .B2 (slo__sro_n134));
NAND2_X1 CLOCK_slo__sro_c990 (.ZN (CLOCK_slo__sro_n1210), .A1 (p_0[4]), .A2 (Multiplier[4]));
XNOR2_X2 slo__sro_c77 (.ZN (p_1[28]), .A (CLOCK_slo__mro_n1162), .B (n_28));
NAND2_X1 slo__sro_c104 (.ZN (slo__sro_n170), .A1 (p_0[29]), .A2 (Multiplier[29]));
NOR2_X1 slo__sro_c105 (.ZN (slo__sro_n169), .A1 (p_0[29]), .A2 (Multiplier[29]));
OAI21_X1 slo__sro_c106 (.ZN (n_30), .A (slo__sro_n170), .B1 (slo__sro_n171), .B2 (slo__sro_n169));
XNOR2_X1 slo__sro_c107 (.ZN (slo__sro_n168), .A (p_0[29]), .B (Multiplier[29]));
XNOR2_X2 slo__sro_c108 (.ZN (p_1[29]), .A (slo__sro_n168), .B (slo__sro_n133));
NAND2_X1 slo__sro_c146 (.ZN (slo__sro_n215), .A1 (n_14), .A2 (Multiplier[14]));
NOR2_X1 slo__sro_c147 (.ZN (slo__sro_n214), .A1 (n_14), .A2 (Multiplier[14]));
OAI21_X2 slo__sro_c148 (.ZN (n_15), .A (slo__sro_n215), .B1 (slo__sro_n214), .B2 (slo__sro_n216));
XNOR2_X1 slo__sro_c149 (.ZN (slo__sro_n213), .A (n_14), .B (Multiplier[14]));
XNOR2_X1 slo__sro_c150 (.ZN (p_1[14]), .A (slo__sro_n213), .B (p_0[14]));
OAI21_X1 slo__sro_c186 (.ZN (slo__sro_n256), .A (p_0[15]), .B1 (n_15), .B2 (Multiplier[15]));
NAND2_X1 slo__sro_c187 (.ZN (n_16), .A1 (slo__sro_n256), .A2 (slo__sro_n257));
XNOR2_X1 slo__sro_c188 (.ZN (slo__sro_n255), .A (n_15), .B (Multiplier[15]));
XNOR2_X1 slo__sro_c189 (.ZN (p_1[15]), .A (slo__sro_n255), .B (p_0[15]));
NAND2_X1 slo__sro_c198 (.ZN (slo__sro_n271), .A1 (p_0[10]), .A2 (Multiplier[10]));
NOR2_X1 slo__sro_c199 (.ZN (slo__sro_n270), .A1 (p_0[10]), .A2 (Multiplier[10]));
OAI21_X1 slo__sro_c200 (.ZN (slo__sro_n269), .A (slo__sro_n271), .B1 (slo__sro_n272), .B2 (slo__sro_n270));
XNOR2_X1 slo__sro_c201 (.ZN (slo__sro_n268), .A (p_0[10]), .B (Multiplier[10]));
XNOR2_X1 slo__sro_c202 (.ZN (p_1[10]), .A (slo__sro_n268), .B (n_10));
NAND2_X1 slo__sro_c326 (.ZN (slo__sro_n447), .A1 (p_0[17]), .A2 (Multiplier[17]));
NOR2_X2 slo__sro_c327 (.ZN (slo__sro_n446), .A1 (p_0[17]), .A2 (Multiplier[17]));
OAI21_X2 slo__sro_c328 (.ZN (n_18), .A (slo__sro_n447), .B1 (slo__n843), .B2 (slo__sro_n446));
XNOR2_X1 slo__sro_c329 (.ZN (slo__sro_n445), .A (p_0[17]), .B (Multiplier[17]));
XNOR2_X1 slo__sro_c330 (.ZN (p_1[17]), .A (slo__sro_n445), .B (n_17));
NAND2_X1 slo__sro_c526 (.ZN (slo__sro_n660), .A1 (n_21), .A2 (Multiplier[21]));
NOR2_X1 slo__sro_c527 (.ZN (slo__sro_n659), .A1 (n_21), .A2 (Multiplier[21]));
OAI21_X1 slo__sro_c528 (.ZN (n_22), .A (slo__sro_n660), .B1 (slo__sro_n659), .B2 (slo__sro_n661));
XNOR2_X1 slo__sro_c529 (.ZN (slo__sro_n658), .A (n_21), .B (Multiplier[21]));
XNOR2_X1 slo__sro_c530 (.ZN (p_1[21]), .A (slo__sro_n658), .B (p_0[21]));
NAND2_X1 slo__sro_c590 (.ZN (slo__sro_n767), .A1 (p_0[12]), .A2 (Multiplier[12]));
NOR2_X1 slo__sro_c591 (.ZN (slo__sro_n766), .A1 (p_0[12]), .A2 (Multiplier[12]));
OAI21_X1 slo__sro_c592 (.ZN (n_13), .A (slo__sro_n767), .B1 (slo__sro_n768), .B2 (slo__sro_n766));
XNOR2_X1 slo__sro_c593 (.ZN (slo__sro_n765), .A (p_0[12]), .B (Multiplier[12]));
XNOR2_X1 slo__sro_c594 (.ZN (p_1[12]), .A (slo__sro_n765), .B (n_12));
XNOR2_X1 slo__mro_c610 (.ZN (p_1[19]), .A (slo__mro_n786), .B (p_0[19]));
NAND2_X1 slo__sro_c638 (.ZN (slo__sro_n828), .A1 (p_0[18]), .A2 (Multiplier[18]));
NAND2_X2 slo__sro_c639 (.ZN (slo__sro_n827), .A1 (n_18), .A2 (Multiplier[18]));
NAND2_X2 slo__sro_c640 (.ZN (slo__sro_n826), .A1 (n_18), .A2 (p_0[18]));
NAND3_X2 slo__sro_c641 (.ZN (n_19), .A1 (slo__sro_n827), .A2 (slo__sro_n826), .A3 (slo__sro_n828));
XNOR2_X1 slo__sro_c642 (.ZN (slo__sro_n825), .A (p_0[18]), .B (Multiplier[18]));
XNOR2_X1 slo__sro_c643 (.ZN (p_1[18]), .A (slo__sro_n825), .B (n_18));
INV_X1 CLOCK_slo__sro_c843 (.ZN (CLOCK_slo__sro_n1068), .A (n_23));
NOR2_X1 CLOCK_slo__sro_c845 (.ZN (CLOCK_slo__sro_n1066), .A1 (p_0[23]), .A2 (Multiplier[23]));
OAI21_X2 CLOCK_slo__sro_c846 (.ZN (CLOCK_slo__sro_n1065), .A (CLOCK_slo__sro_n1067)
    , .B1 (CLOCK_slo__sro_n1068), .B2 (CLOCK_slo__sro_n1066));
XNOR2_X1 CLOCK_slo__sro_c847 (.ZN (CLOCK_slo__sro_n1064), .A (p_0[23]), .B (Multiplier[23]));
XNOR2_X1 CLOCK_slo__sro_c848 (.ZN (p_1[23]), .A (CLOCK_slo__sro_n1064), .B (n_23));
XNOR2_X1 CLOCK_slo__mro_c858 (.ZN (p_1[24]), .A (CLOCK_slo__mro_n1081), .B (p_0[24]));
NOR2_X1 CLOCK_slo__sro_c878 (.ZN (CLOCK_slo__sro_n1101), .A1 (p_0[16]), .A2 (Multiplier[16]));
OAI21_X2 CLOCK_slo__sro_c879 (.ZN (n_17), .A (CLOCK_slo__sro_n1102), .B1 (CLOCK_slo__sro_n1103), .B2 (CLOCK_slo__sro_n1101));
XNOR2_X1 CLOCK_slo__sro_c880 (.ZN (CLOCK_slo__sro_n1100), .A (p_0[16]), .B (Multiplier[16]));
XNOR2_X1 CLOCK_slo__sro_c881 (.ZN (p_1[16]), .A (CLOCK_slo__sro_n1100), .B (n_16));
NAND2_X1 CLOCK_slo__sro_c991 (.ZN (CLOCK_slo__sro_n1209), .A1 (n_4), .A2 (Multiplier[4]));
NAND2_X1 CLOCK_slo__sro_c992 (.ZN (CLOCK_slo__sro_n1208), .A1 (p_0[4]), .A2 (n_4));
NAND3_X1 CLOCK_slo__sro_c993 (.ZN (CLOCK_slo__sro_n1207), .A1 (CLOCK_slo__sro_n1208)
    , .A2 (CLOCK_slo__sro_n1210), .A3 (CLOCK_slo__sro_n1209));
XNOR2_X1 CLOCK_slo__sro_c994 (.ZN (CLOCK_slo__sro_n1206), .A (p_0[4]), .B (Multiplier[4]));
XNOR2_X1 CLOCK_slo__sro_c995 (.ZN (p_1[4]), .A (CLOCK_slo__sro_n1206), .B (n_4));
NAND2_X1 CLOCK_slo__sro_c1016 (.ZN (CLOCK_slo__sro_n1235), .A1 (p_0[8]), .A2 (Multiplier[8]));
NOR2_X1 CLOCK_slo__sro_c1017 (.ZN (CLOCK_slo__sro_n1234), .A1 (p_0[8]), .A2 (Multiplier[8]));
OAI21_X1 CLOCK_slo__sro_c1018 (.ZN (n_9), .A (CLOCK_slo__sro_n1235), .B1 (CLOCK_slo__sro_n1236), .B2 (CLOCK_slo__sro_n1234));
XNOR2_X1 CLOCK_slo__sro_c1019 (.ZN (CLOCK_slo__sro_n1233), .A (p_0[8]), .B (Multiplier[8]));
XNOR2_X1 CLOCK_slo__sro_c1020 (.ZN (p_1[8]), .A (CLOCK_slo__sro_n1233), .B (n_8));
NOR2_X1 CLOCK_slo__sro_c1387 (.ZN (CLOCK_slo__sro_n1598), .A1 (p_0[11]), .A2 (Multiplier[11]));
INV_X1 CLOCK_slo__sro_c1227 (.ZN (CLOCK_slo__sro_n1452), .A (n_27));
NAND2_X1 CLOCK_slo__sro_c1228 (.ZN (CLOCK_slo__sro_n1451), .A1 (p_0[27]), .A2 (Multiplier[27]));
NOR2_X1 CLOCK_slo__sro_c1229 (.ZN (CLOCK_slo__sro_n1450), .A1 (p_0[27]), .A2 (Multiplier[27]));
OAI21_X4 CLOCK_slo__sro_c1083 (.ZN (n_14), .A (slo__sro_n61), .B1 (slo__sro_n62), .B2 (slo__sro_n60));
XNOR2_X1 CLOCK_slo__sro_c1231 (.ZN (CLOCK_slo__sro_n1449), .A (p_0[27]), .B (Multiplier[27]));
XNOR2_X1 CLOCK_slo__sro_c1232 (.ZN (p_1[27]), .A (CLOCK_slo__sro_n1449), .B (n_27));
XNOR2_X1 CLOCK_slo__sro_c1390 (.ZN (p_1[11]), .A (slo__sro_n269), .B (CLOCK_slo__sro_n1597));

endmodule //datapath__0_161

module datapath__0_157 (p_0, p_1, p_2);

output [31:0] p_2;
input [31:0] p_0;
input [31:0] p_1;
wire slo__sro_n529;
wire slo__sro_n437;
wire n_1;
wire n_3;
wire n_4;
wire n_5;
wire n_6;
wire n_7;
wire n_8;
wire n_10;
wire n_12;
wire n_14;
wire n_15;
wire n_16;
wire slo__sro_n312;
wire n_19;
wire slo__sro_n341;
wire n_21;
wire n_22;
wire n_23;
wire CLOCK_slo__sro_n1406;
wire n_27;
wire CLOCK_slo__sro_n1345;
wire n_29;
wire n_30;
wire n_32;
wire n_0;
wire n_34;
wire n_33;
wire n_31;
wire slo__sro_n134;
wire slo__sro_n135;
wire slo__sro_n136;
wire slo__sro_n137;
wire slo__sro_n138;
wire slo__sro_n308;
wire slo__sro_n309;
wire slo__sro_n310;
wire slo__sro_n311;
wire slo__sro_n102;
wire slo__sro_n103;
wire slo__sro_n104;
wire slo__sro_n105;
wire slo__sro_n106;
wire slo__sro_n177;
wire slo__sro_n178;
wire slo__sro_n179;
wire slo__sro_n180;
wire slo__sro_n325;
wire slo__sro_n326;
wire slo__sro_n327;
wire slo__sro_n328;
wire slo__sro_n264;
wire slo__sro_n265;
wire slo__sro_n266;
wire slo__sro_n267;
wire slo__sro_n268;
wire slo__sro_n342;
wire slo__sro_n343;
wire slo__sro_n420;
wire slo__sro_n421;
wire slo__sro_n422;
wire slo__sro_n423;
wire slo__sro_n514;
wire slo__sro_n515;
wire slo__sro_n516;
wire slo__sro_n517;
wire slo__sro_n530;
wire slo__sro_n531;
wire slo__sro_n532;
wire slo__sro_n747;
wire slo__sro_n748;
wire slo__sro_n749;
wire slo__sro_n750;
wire slo__sro_n798;
wire slo__sro_n799;
wire slo__sro_n800;
wire slo__sro_n801;
wire slo__sro_n855;
wire slo__sro_n856;
wire slo__sro_n857;
wire slo__sro_n858;
wire slo__sro_n883;
wire slo__sro_n884;
wire slo__sro_n885;
wire slo__sro_n886;
wire slo__sro_n887;
wire slo__sro_n915;
wire slo__sro_n916;
wire slo__sro_n917;
wire slo__sro_n918;
wire CLOCK_slo__sro_n1405;
wire slo__n1123;
wire CLOCK_slo__sro_n1285;
wire CLOCK_slo__sro_n1286;
wire CLOCK_slo__sro_n1287;
wire CLOCK_slo__sro_n1288;
wire CLOCK_slo__sro_n1308;
wire CLOCK_slo__sro_n1309;
wire CLOCK_slo__sro_n1310;
wire CLOCK_slo__mro_n1324;
wire CLOCK_slo__sro_n1346;
wire CLOCK_slo__sro_n1347;
wire CLOCK_slo__sro_n1348;
wire CLOCK_slo__sro_n1349;
wire CLOCK_slo__sro_n1407;
wire CLOCK_slo__sro_n1408;


INV_X1 i_36 (.ZN (n_34), .A (p_0[30]));
INV_X1 i_35 (.ZN (n_33), .A (p_1[30]));
INV_X1 i_34 (.ZN (n_32), .A (n_30));
XOR2_X1 i_32 (.Z (p_2[31]), .A (p_0[31]), .B (n_31));
OAI22_X1 i_31 (.ZN (n_0), .A1 (n_34), .A2 (p_1[30]), .B1 (p_0[30]), .B2 (n_33));
XNOR2_X1 i_0 (.ZN (p_2[30]), .A (n_32), .B (n_0));
FA_X1 i_30 (.CO (n_30), .S (p_2[29]), .A (p_0[29]), .B (p_1[29]), .CI (n_29));
FA_X1 i_29 (.CO (n_29), .S (p_2[28]), .A (p_0[28]), .B (p_1[28]), .CI (slo__sro_n326));
INV_X1 slo__sro_c256 (.ZN (slo__sro_n343), .A (n_4));
FA_X1 i_27 (.CO (n_27), .S (p_2[26]), .A (p_0[26]), .B (p_1[26]), .CI (slo__sro_n748));
INV_X1 slo__sro_c535 (.ZN (slo__sro_n801), .A (n_3));
NOR2_X1 CLOCK_slo__sro_c918 (.ZN (CLOCK_slo__sro_n1407), .A1 (n_33), .A2 (p_0[30]));
NAND2_X1 slo__sro_c108 (.ZN (slo__sro_n179), .A1 (p_1[17]), .A2 (p_0[17]));
FA_X1 i_23 (.CO (n_23), .S (p_2[22]), .A (p_0[22]), .B (p_1[22]), .CI (n_22));
FA_X1 i_22 (.CO (n_22), .S (p_2[21]), .A (p_0[21]), .B (p_1[21]), .CI (n_21));
FA_X1 i_21 (.CO (n_21), .S (p_2[20]), .A (p_0[20]), .B (p_1[20]), .CI (slo__sro_n265));
OAI21_X1 slo__sro_c259 (.ZN (n_5), .A (slo__sro_n342), .B1 (slo__sro_n343), .B2 (slo__sro_n341));
NAND2_X1 slo__sro_c379 (.ZN (slo__sro_n532), .A1 (p_1[10]), .A2 (p_0[10]));
OAI21_X1 slo__sro_c245 (.ZN (slo__sro_n327), .A (n_27), .B1 (p_1[27]), .B2 (p_0[27]));
INV_X1 slo__sro_c623 (.ZN (slo__sro_n918), .A (CLOCK_slo__sro_n1286));
FA_X1 i_16 (.CO (n_16), .S (p_2[15]), .A (p_0[15]), .B (p_1[15]), .CI (n_15));
FA_X1 i_15 (.CO (n_15), .S (p_2[14]), .A (p_0[14]), .B (p_1[14]), .CI (n_14));
INV_X1 CLOCK_slo__sro_c917 (.ZN (CLOCK_slo__sro_n1408), .A (n_30));
NAND2_X1 CLOCK_slo__sro_c824 (.ZN (CLOCK_slo__sro_n1310), .A1 (p_1[11]), .A2 (p_0[11]));
XNOR2_X1 CLOCK_slo__mro_c839 (.ZN (CLOCK_slo__mro_n1324), .A (n_4), .B (p_0[4]));
NAND2_X1 slo__sro_c511 (.ZN (slo__sro_n750), .A1 (p_1[25]), .A2 (p_0[25]));
FA_X1 i_10 (.CO (n_10), .S (p_2[9]), .A (p_0[9]), .B (p_1[9]), .CI (slo__sro_n309));
NAND2_X1 slo__sro_c244 (.ZN (slo__sro_n328), .A1 (p_1[27]), .A2 (p_0[27]));
XNOR2_X1 slo__sro_c324 (.ZN (slo__sro_n437), .A (p_1[17]), .B (p_0[17]));
FA_X1 i_7 (.CO (n_7), .S (p_2[6]), .A (p_0[6]), .B (p_1[6]), .CI (n_6));
FA_X1 i_6 (.CO (n_6), .S (p_2[5]), .A (p_0[5]), .B (p_1[5]), .CI (n_5));
NAND2_X1 CLOCK_slo__sro_c806 (.ZN (CLOCK_slo__sro_n1288), .A1 (p_1[12]), .A2 (p_0[12]));
INV_X1 slo__sro_c576 (.ZN (slo__sro_n858), .A (p_1[2]));
INV_X1 slo__sro_c596 (.ZN (slo__sro_n887), .A (n_16));
INV_X1 slo__sro_c230 (.ZN (slo__sro_n312), .A (n_8));
HA_X1 i_1 (.CO (n_1), .S (p_2[0]), .A (p_0[0]), .B (p_1[0]));
INV_X2 slo__sro_c67 (.ZN (slo__sro_n138), .A (p_1[1]));
NAND2_X1 slo__sro_c68 (.ZN (slo__sro_n137), .A1 (n_1), .A2 (p_0[1]));
NOR2_X1 slo__sro_c69 (.ZN (slo__sro_n136), .A1 (n_1), .A2 (p_0[1]));
OAI21_X2 slo__sro_c70 (.ZN (slo__sro_n135), .A (slo__sro_n137), .B1 (slo__sro_n138), .B2 (slo__sro_n136));
XNOR2_X2 slo__sro_c71 (.ZN (slo__sro_n134), .A (n_1), .B (p_0[1]));
XNOR2_X1 slo__sro_c72 (.ZN (p_2[1]), .A (p_1[1]), .B (slo__sro_n134));
NAND2_X1 slo__sro_c231 (.ZN (slo__sro_n311), .A1 (p_1[8]), .A2 (p_0[8]));
NOR2_X1 slo__sro_c232 (.ZN (slo__sro_n310), .A1 (p_1[8]), .A2 (p_0[8]));
OAI21_X1 slo__sro_c233 (.ZN (slo__sro_n309), .A (slo__sro_n311), .B1 (slo__sro_n312), .B2 (slo__sro_n310));
XNOR2_X1 slo__sro_c234 (.ZN (slo__sro_n308), .A (p_1[8]), .B (p_0[8]));
XNOR2_X1 slo__sro_c235 (.ZN (p_2[8]), .A (slo__sro_n308), .B (n_8));
INV_X1 slo__sro_c107 (.ZN (slo__sro_n180), .A (slo__sro_n884));
INV_X1 slo__sro_c40 (.ZN (slo__sro_n106), .A (n_23));
NAND2_X1 slo__sro_c41 (.ZN (slo__sro_n105), .A1 (p_1[23]), .A2 (p_0[23]));
NOR2_X1 slo__sro_c42 (.ZN (slo__sro_n104), .A1 (p_1[23]), .A2 (p_0[23]));
OAI21_X1 slo__sro_c43 (.ZN (slo__sro_n103), .A (slo__sro_n105), .B1 (slo__sro_n106), .B2 (slo__sro_n104));
XNOR2_X1 slo__sro_c44 (.ZN (slo__sro_n102), .A (p_1[23]), .B (p_0[23]));
XNOR2_X1 slo__sro_c45 (.ZN (p_2[23]), .A (slo__sro_n102), .B (n_23));
NOR2_X1 slo__sro_c109 (.ZN (slo__sro_n178), .A1 (p_1[17]), .A2 (p_0[17]));
OAI21_X1 slo__sro_c110 (.ZN (slo__sro_n177), .A (slo__sro_n179), .B1 (slo__sro_n180), .B2 (slo__sro_n178));
INV_X1 slo__sro_c364 (.ZN (slo__sro_n517), .A (slo__sro_n177));
INV_X1 slo__sro_c308 (.ZN (slo__sro_n423), .A (n_7));
NAND2_X1 slo__sro_c246 (.ZN (slo__sro_n326), .A1 (slo__sro_n328), .A2 (slo__sro_n327));
XNOR2_X1 slo__sro_c247 (.ZN (slo__sro_n325), .A (p_1[27]), .B (p_0[27]));
XNOR2_X1 slo__sro_c248 (.ZN (p_2[27]), .A (slo__sro_n325), .B (n_27));
NAND2_X1 slo__sro_c257 (.ZN (slo__sro_n342), .A1 (p_1[4]), .A2 (p_0[4]));
NOR2_X1 slo__sro_c258 (.ZN (slo__sro_n341), .A1 (p_1[4]), .A2 (p_0[4]));
INV_X1 slo__sro_c190 (.ZN (slo__sro_n268), .A (n_19));
NAND2_X1 slo__sro_c191 (.ZN (slo__sro_n267), .A1 (p_1[19]), .A2 (p_0[19]));
NOR2_X1 slo__sro_c192 (.ZN (slo__sro_n266), .A1 (p_1[19]), .A2 (p_0[19]));
OAI21_X1 slo__sro_c193 (.ZN (slo__sro_n265), .A (slo__sro_n267), .B1 (slo__sro_n268), .B2 (slo__sro_n266));
XNOR2_X1 slo__sro_c194 (.ZN (slo__sro_n264), .A (p_1[19]), .B (p_0[19]));
XNOR2_X1 slo__sro_c195 (.ZN (p_2[19]), .A (slo__sro_n264), .B (n_19));
INV_X1 CLOCK_slo__sro_c858 (.ZN (CLOCK_slo__sro_n1349), .A (slo__sro_n103));
NAND2_X1 CLOCK_slo__sro_c859 (.ZN (CLOCK_slo__sro_n1348), .A1 (p_1[24]), .A2 (p_0[24]));
XNOR2_X1 slo__sro_c300 (.ZN (p_2[17]), .A (slo__sro_n437), .B (slo__sro_n884));
NAND2_X1 slo__sro_c309 (.ZN (slo__sro_n422), .A1 (p_1[7]), .A2 (p_0[7]));
NOR2_X1 slo__sro_c310 (.ZN (slo__sro_n421), .A1 (p_1[7]), .A2 (p_0[7]));
OAI21_X1 slo__sro_c311 (.ZN (n_8), .A (slo__sro_n422), .B1 (slo__sro_n423), .B2 (slo__sro_n421));
XNOR2_X1 slo__sro_c312 (.ZN (slo__sro_n420), .A (p_1[7]), .B (p_0[7]));
XNOR2_X1 slo__sro_c313 (.ZN (p_2[7]), .A (slo__sro_n420), .B (n_7));
NAND2_X1 slo__sro_c365 (.ZN (slo__sro_n516), .A1 (p_1[18]), .A2 (p_0[18]));
NOR2_X1 slo__sro_c366 (.ZN (slo__sro_n515), .A1 (p_1[18]), .A2 (p_0[18]));
OAI21_X1 slo__sro_c367 (.ZN (n_19), .A (slo__sro_n516), .B1 (slo__sro_n517), .B2 (slo__sro_n515));
XNOR2_X2 slo__sro_c368 (.ZN (slo__sro_n514), .A (p_1[18]), .B (p_0[18]));
XNOR2_X1 slo__sro_c369 (.ZN (p_2[18]), .A (slo__sro_n514), .B (slo__sro_n177));
NOR2_X1 slo__sro_c380 (.ZN (slo__sro_n531), .A1 (p_1[10]), .A2 (p_0[10]));
OAI21_X1 slo__sro_c381 (.ZN (slo__sro_n530), .A (slo__sro_n532), .B1 (slo__sro_n531), .B2 (slo__n1123));
XNOR2_X1 slo__sro_c382 (.ZN (slo__sro_n529), .A (p_1[10]), .B (p_0[10]));
XNOR2_X1 slo__sro_c383 (.ZN (p_2[10]), .A (slo__sro_n529), .B (n_10));
OAI21_X1 slo__sro_c512 (.ZN (slo__sro_n749), .A (CLOCK_slo__sro_n1346), .B1 (p_1[25]), .B2 (p_0[25]));
NAND2_X1 slo__sro_c513 (.ZN (slo__sro_n748), .A1 (slo__sro_n749), .A2 (slo__sro_n750));
XNOR2_X1 slo__sro_c514 (.ZN (slo__sro_n747), .A (p_1[25]), .B (p_0[25]));
XNOR2_X1 slo__sro_c515 (.ZN (p_2[25]), .A (slo__sro_n747), .B (CLOCK_slo__sro_n1346));
NAND2_X1 slo__sro_c536 (.ZN (slo__sro_n800), .A1 (p_1[3]), .A2 (p_0[3]));
NOR2_X1 slo__sro_c537 (.ZN (slo__sro_n799), .A1 (p_1[3]), .A2 (p_0[3]));
OAI21_X1 slo__sro_c538 (.ZN (n_4), .A (slo__sro_n800), .B1 (slo__sro_n799), .B2 (slo__sro_n801));
XNOR2_X2 slo__sro_c539 (.ZN (slo__sro_n798), .A (p_1[3]), .B (p_0[3]));
XNOR2_X1 slo__sro_c540 (.ZN (p_2[3]), .A (slo__sro_n798), .B (n_3));
NAND2_X1 slo__sro_c577 (.ZN (slo__sro_n857), .A1 (slo__sro_n135), .A2 (p_0[2]));
NOR2_X1 slo__sro_c578 (.ZN (slo__sro_n856), .A1 (slo__sro_n135), .A2 (p_0[2]));
OAI21_X2 slo__sro_c579 (.ZN (n_3), .A (slo__sro_n857), .B1 (slo__sro_n858), .B2 (slo__sro_n856));
XNOR2_X2 slo__sro_c580 (.ZN (slo__sro_n855), .A (slo__sro_n135), .B (p_0[2]));
XNOR2_X2 slo__sro_c581 (.ZN (p_2[2]), .A (slo__sro_n855), .B (p_1[2]));
NAND2_X1 slo__sro_c597 (.ZN (slo__sro_n886), .A1 (p_1[16]), .A2 (p_0[16]));
NOR2_X1 slo__sro_c598 (.ZN (slo__sro_n885), .A1 (p_1[16]), .A2 (p_0[16]));
OAI21_X1 slo__sro_c599 (.ZN (slo__sro_n884), .A (slo__sro_n886), .B1 (slo__sro_n887), .B2 (slo__sro_n885));
XNOR2_X1 slo__sro_c600 (.ZN (slo__sro_n883), .A (p_1[16]), .B (p_0[16]));
XNOR2_X1 slo__sro_c601 (.ZN (p_2[16]), .A (slo__sro_n883), .B (n_16));
NAND2_X1 slo__sro_c624 (.ZN (slo__sro_n917), .A1 (p_1[13]), .A2 (p_0[13]));
NOR2_X1 slo__sro_c625 (.ZN (slo__sro_n916), .A1 (p_1[13]), .A2 (p_0[13]));
OAI21_X1 slo__sro_c626 (.ZN (n_14), .A (slo__sro_n917), .B1 (slo__sro_n916), .B2 (slo__sro_n918));
XNOR2_X1 slo__sro_c627 (.ZN (slo__sro_n915), .A (p_1[13]), .B (p_0[13]));
XNOR2_X1 slo__sro_c628 (.ZN (p_2[13]), .A (slo__sro_n915), .B (CLOCK_slo__sro_n1286));
INV_X1 slo__L1_c740 (.ZN (slo__n1123), .A (n_10));
OAI21_X1 CLOCK_slo__sro_c807 (.ZN (CLOCK_slo__sro_n1287), .A (n_12), .B1 (p_1[12]), .B2 (p_0[12]));
NAND2_X1 CLOCK_slo__sro_c808 (.ZN (CLOCK_slo__sro_n1286), .A1 (CLOCK_slo__sro_n1287), .A2 (CLOCK_slo__sro_n1288));
XNOR2_X1 CLOCK_slo__sro_c809 (.ZN (CLOCK_slo__sro_n1285), .A (p_1[12]), .B (p_0[12]));
XNOR2_X1 CLOCK_slo__sro_c810 (.ZN (p_2[12]), .A (CLOCK_slo__sro_n1285), .B (n_12));
OAI21_X1 CLOCK_slo__sro_c825 (.ZN (CLOCK_slo__sro_n1309), .A (slo__sro_n530), .B1 (p_1[11]), .B2 (p_0[11]));
NAND2_X1 CLOCK_slo__sro_c826 (.ZN (n_12), .A1 (CLOCK_slo__sro_n1309), .A2 (CLOCK_slo__sro_n1310));
XNOR2_X1 CLOCK_slo__sro_c827 (.ZN (CLOCK_slo__sro_n1308), .A (slo__sro_n530), .B (p_0[11]));
XNOR2_X1 CLOCK_slo__sro_c828 (.ZN (p_2[11]), .A (CLOCK_slo__sro_n1308), .B (p_1[11]));
XNOR2_X1 CLOCK_slo__mro_c840 (.ZN (p_2[4]), .A (CLOCK_slo__mro_n1324), .B (p_1[4]));
NOR2_X1 CLOCK_slo__sro_c860 (.ZN (CLOCK_slo__sro_n1347), .A1 (p_1[24]), .A2 (p_0[24]));
OAI21_X1 CLOCK_slo__sro_c861 (.ZN (CLOCK_slo__sro_n1346), .A (CLOCK_slo__sro_n1348)
    , .B1 (CLOCK_slo__sro_n1349), .B2 (CLOCK_slo__sro_n1347));
XNOR2_X1 CLOCK_slo__sro_c862 (.ZN (CLOCK_slo__sro_n1345), .A (p_1[24]), .B (p_0[24]));
XNOR2_X1 CLOCK_slo__sro_c863 (.ZN (p_2[24]), .A (CLOCK_slo__sro_n1345), .B (slo__sro_n103));
NAND2_X1 CLOCK_slo__sro_c919 (.ZN (CLOCK_slo__sro_n1406), .A1 (CLOCK_slo__sro_n1408), .A2 (CLOCK_slo__sro_n1407));
OR2_X1 CLOCK_slo__sro_c920 (.ZN (CLOCK_slo__sro_n1405), .A1 (p_1[30]), .A2 (n_34));
OAI21_X1 CLOCK_slo__sro_c921 (.ZN (n_31), .A (CLOCK_slo__sro_n1406), .B1 (n_32), .B2 (CLOCK_slo__sro_n1405));

endmodule //datapath__0_157

module datapath__0_156 (Multiplier, p_0, p_1);

output [31:0] p_1;
input [31:0] Multiplier;
input [31:0] p_0;
wire n_1;
wire n_2;
wire n_3;
wire n_4;
wire n_5;
wire n_6;
wire n_7;
wire slo__sro_n729;
wire CLOCK_slo__sro_n1418;
wire n_11;
wire n_12;
wire n_13;
wire CLOCK_slo__sro_n1108;
wire n_15;
wire slo__sro_n361;
wire n_18;
wire n_19;
wire slo__sro_n487;
wire CLOCK_slo__sro_n1107;
wire n_22;
wire n_23;
wire n_24;
wire n_25;
wire n_26;
wire n_28;
wire n_29;
wire n_30;
wire n_32;
wire n_0;
wire n_34;
wire n_33;
wire n_31;
wire slo__sro_n59;
wire slo__sro_n60;
wire slo__sro_n61;
wire slo__sro_n62;
wire slo__sro_n63;
wire slo__sro_n77;
wire slo__sro_n78;
wire slo__sro_n79;
wire slo__sro_n730;
wire slo__sro_n106;
wire slo__sro_n107;
wire slo__sro_n108;
wire slo__sro_n109;
wire slo__sro_n146;
wire slo__sro_n147;
wire slo__sro_n148;
wire slo__sro_n149;
wire slo__sro_n161;
wire slo__sro_n163;
wire slo__sro_n357;
wire slo__sro_n358;
wire slo__sro_n359;
wire slo__sro_n360;
wire slo__sro_n189;
wire slo__sro_n190;
wire slo__sro_n191;
wire slo__sro_n192;
wire slo__sro_n193;
wire slo__sro_n488;
wire slo__sro_n489;
wire slo__sro_n490;
wire slo__sro_n491;
wire slo__xsl_n643;
wire slo__sro_n247;
wire slo__sro_n248;
wire slo__sro_n249;
wire slo__sro_n250;
wire slo__sro_n251;
wire slo__sro_n731;
wire slo__sro_n732;
wire slo__sro_n733;
wire CLOCK_slo__mro_n1025;
wire slo__sro_n464;
wire slo__sro_n465;
wire slo__sro_n466;
wire slo__sro_n467;
wire slo__sro_n468;
wire CLOCK_slo__sro_n1109;
wire CLOCK_slo__sro_n1110;
wire CLOCK_slo__sro_n1135;
wire CLOCK_slo__sro_n1136;
wire CLOCK_slo__sro_n1137;
wire CLOCK_slo__sro_n1138;
wire CLOCK_slo__sro_n1184;
wire CLOCK_slo__sro_n1185;
wire CLOCK_slo__sro_n1186;
wire CLOCK_slo__sro_n1187;
wire CLOCK_slo__sro_n1188;
wire CLOCK_slo__sro_n1417;
wire CLOCK_slo__sro_n1419;
wire slo__sro_n861;
wire slo__sro_n862;
wire slo__sro_n863;
wire slo__sro_n864;


INV_X1 i_36 (.ZN (n_34), .A (Multiplier[30]));
INV_X1 i_35 (.ZN (n_33), .A (p_0[30]));
INV_X1 i_34 (.ZN (n_32), .A (n_30));
OAI33_X1 i_33 (.ZN (n_31), .A1 (n_34), .A2 (p_0[30]), .A3 (n_32), .B1 (n_30), .B2 (n_33), .B3 (Multiplier[30]));
XOR2_X1 i_32 (.Z (p_1[31]), .A (Multiplier[31]), .B (n_31));
OAI22_X1 i_31 (.ZN (n_0), .A1 (n_34), .A2 (p_0[30]), .B1 (Multiplier[30]), .B2 (n_33));
XNOR2_X1 i_0 (.ZN (p_1[30]), .A (n_32), .B (n_0));
FA_X1 i_30 (.CO (n_30), .S (p_1[29]), .A (Multiplier[29]), .B (p_0[29]), .CI (n_29));
NAND2_X1 CLOCK_slo__sro_c918 (.ZN (CLOCK_slo__sro_n1188), .A1 (p_0[9]), .A2 (Multiplier[9]));
NAND2_X1 slo__sro_c98 (.ZN (slo__sro_n163), .A1 (p_0[25]), .A2 (Multiplier[25]));
INV_X1 slo__sro_c42 (.ZN (slo__sro_n109), .A (n_23));
INV_X1 slo__sro_c333 (.ZN (slo__sro_n491), .A (n_7));
FA_X1 i_25 (.CO (n_25), .S (p_1[24]), .A (Multiplier[24]), .B (p_0[24]), .CI (n_24));
NAND2_X1 slo__sro_c82 (.ZN (slo__sro_n149), .A1 (p_0[27]), .A2 (Multiplier[27]));
FA_X1 i_23 (.CO (n_23), .S (p_1[22]), .A (Multiplier[22]), .B (p_0[22]), .CI (n_22));
FA_X1 i_22 (.CO (n_22), .S (p_1[21]), .A (Multiplier[21]), .B (p_0[21]), .CI (slo__sro_n60));
OAI21_X1 slo__sro_c548 (.ZN (slo__sro_n730), .A (slo__sro_n732), .B1 (slo__sro_n731), .B2 (slo__sro_n733));
NAND2_X1 slo__sro_c334 (.ZN (slo__sro_n490), .A1 (p_0[7]), .A2 (Multiplier[7]));
FA_X1 i_19 (.CO (n_19), .S (p_1[18]), .A (Multiplier[18]), .B (p_0[18]), .CI (n_18));
FA_X1 i_18 (.CO (n_18), .S (p_1[17]), .A (Multiplier[17]), .B (p_0[17]), .CI (slo__sro_n730));
XNOR2_X2 CLOCK_slo__mro_c765 (.ZN (CLOCK_slo__mro_n1025), .A (p_0[26]), .B (Multiplier[26]));
XNOR2_X1 slo__sro_c237 (.ZN (p_1[19]), .A (slo__sro_n357), .B (n_19));
FA_X1 i_15 (.CO (n_15), .S (p_1[14]), .A (Multiplier[14]), .B (p_0[14]), .CI (slo__sro_n465));
OAI21_X1 CLOCK_slo__sro_c844 (.ZN (n_2), .A (CLOCK_slo__sro_n1109), .B1 (CLOCK_slo__sro_n1110), .B2 (CLOCK_slo__sro_n1108));
FA_X1 i_13 (.CO (n_13), .S (p_1[12]), .A (Multiplier[12]), .B (p_0[12]), .CI (n_12));
FA_X1 i_12 (.CO (n_12), .S (p_1[11]), .A (Multiplier[11]), .B (p_0[11]), .CI (n_11));
NAND2_X1 CLOCK_slo__sro_c1145 (.ZN (CLOCK_slo__sro_n1417), .A1 (n_25), .A2 (CLOCK_slo__sro_n1418));
NOR2_X1 slo__sro_c547 (.ZN (slo__sro_n731), .A1 (slo__sro_n190), .A2 (Multiplier[16]));
INV_X1 slo__sro_c545 (.ZN (slo__sro_n733), .A (p_0[16]));
FA_X1 i_7 (.CO (n_7), .S (p_1[6]), .A (Multiplier[6]), .B (p_0[6]), .CI (n_6));
FA_X1 i_6 (.CO (n_6), .S (p_1[5]), .A (Multiplier[5]), .B (p_0[5]), .CI (n_5));
FA_X1 i_5 (.CO (n_5), .S (p_1[4]), .A (Multiplier[4]), .B (p_0[4]), .CI (n_4));
FA_X1 i_4 (.CO (n_4), .S (p_1[3]), .A (Multiplier[3]), .B (p_0[3]), .CI (n_3));
FA_X1 i_3 (.CO (n_3), .S (p_1[2]), .A (Multiplier[2]), .B (p_0[2]), .CI (n_2));
NAND2_X1 CLOCK_slo__sro_c868 (.ZN (CLOCK_slo__sro_n1138), .A1 (p_0[28]), .A2 (Multiplier[28]));
HA_X1 i_1 (.CO (n_1), .S (p_1[0]), .A (Multiplier[0]), .B (p_0[0]));
INV_X2 slo__sro_c1 (.ZN (slo__sro_n63), .A (slo__sro_n358));
NAND2_X1 slo__sro_c2 (.ZN (slo__sro_n62), .A1 (p_0[20]), .A2 (Multiplier[20]));
NOR2_X1 slo__sro_c3 (.ZN (slo__sro_n61), .A1 (p_0[20]), .A2 (Multiplier[20]));
OAI21_X1 slo__sro_c4 (.ZN (slo__sro_n60), .A (slo__sro_n62), .B1 (slo__sro_n63), .B2 (slo__sro_n61));
XNOR2_X1 slo__sro_c5 (.ZN (slo__sro_n59), .A (p_0[20]), .B (Multiplier[20]));
XNOR2_X1 slo__sro_c6 (.ZN (p_1[20]), .A (slo__sro_n59), .B (slo__sro_n358));
NAND2_X1 slo__sro_c16 (.ZN (slo__sro_n79), .A1 (p_0[26]), .A2 (Multiplier[26]));
NOR2_X2 slo__sro_c17 (.ZN (slo__sro_n78), .A1 (p_0[26]), .A2 (Multiplier[26]));
OAI21_X2 slo__sro_c18 (.ZN (slo__sro_n77), .A (slo__sro_n79), .B1 (slo__sro_n78), .B2 (n_26));
INV_X1 CLOCK_slo__sro_c841 (.ZN (CLOCK_slo__sro_n1110), .A (p_0[1]));
NAND2_X1 CLOCK_slo__sro_c842 (.ZN (CLOCK_slo__sro_n1109), .A1 (n_1), .A2 (Multiplier[1]));
NAND2_X1 slo__sro_c43 (.ZN (slo__sro_n108), .A1 (p_0[23]), .A2 (Multiplier[23]));
NOR2_X1 slo__sro_c44 (.ZN (slo__sro_n107), .A1 (p_0[23]), .A2 (Multiplier[23]));
OAI21_X1 slo__sro_c45 (.ZN (n_24), .A (slo__sro_n108), .B1 (slo__sro_n109), .B2 (slo__sro_n107));
XNOR2_X1 slo__sro_c46 (.ZN (slo__sro_n106), .A (p_0[23]), .B (Multiplier[23]));
XNOR2_X1 slo__sro_c47 (.ZN (p_1[23]), .A (n_23), .B (slo__sro_n106));
NAND2_X1 slo__sro_c83 (.ZN (slo__sro_n148), .A1 (slo__sro_n77), .A2 (Multiplier[27]));
NAND2_X1 slo__sro_c84 (.ZN (slo__sro_n147), .A1 (p_0[27]), .A2 (slo__sro_n77));
NAND3_X1 slo__sro_c85 (.ZN (n_28), .A1 (slo__sro_n149), .A2 (slo__sro_n147), .A3 (slo__sro_n148));
XNOR2_X1 slo__sro_c86 (.ZN (slo__sro_n146), .A (slo__sro_n77), .B (Multiplier[27]));
XNOR2_X1 slo__sro_c87 (.ZN (p_1[27]), .A (slo__sro_n146), .B (p_0[27]));
XNOR2_X2 slo__sro_c549 (.ZN (slo__sro_n729), .A (slo__sro_n190), .B (Multiplier[16]));
XNOR2_X2 slo__sro_c101 (.ZN (slo__sro_n161), .A (p_0[25]), .B (Multiplier[25]));
XNOR2_X1 slo__sro_c102 (.ZN (p_1[25]), .A (slo__sro_n161), .B (n_25));
INV_X1 slo__sro_c232 (.ZN (slo__sro_n361), .A (n_19));
NAND2_X1 slo__sro_c233 (.ZN (slo__sro_n360), .A1 (p_0[19]), .A2 (Multiplier[19]));
NOR2_X1 slo__sro_c234 (.ZN (slo__sro_n359), .A1 (p_0[19]), .A2 (Multiplier[19]));
OAI21_X2 slo__sro_c235 (.ZN (slo__sro_n358), .A (slo__sro_n360), .B1 (slo__sro_n361), .B2 (slo__sro_n359));
XNOR2_X1 slo__sro_c236 (.ZN (slo__sro_n357), .A (p_0[19]), .B (Multiplier[19]));
INV_X2 slo__sro_c123 (.ZN (slo__sro_n193), .A (n_15));
NAND2_X1 slo__sro_c124 (.ZN (slo__sro_n192), .A1 (p_0[15]), .A2 (Multiplier[15]));
NOR2_X2 slo__sro_c125 (.ZN (slo__sro_n191), .A1 (p_0[15]), .A2 (Multiplier[15]));
XNOR2_X2 CLOCK_slo__mro_c766 (.ZN (p_1[26]), .A (CLOCK_slo__mro_n1025), .B (slo__xsl_n643));
XNOR2_X1 slo__sro_c127 (.ZN (slo__sro_n189), .A (p_0[15]), .B (Multiplier[15]));
XNOR2_X1 slo__sro_c128 (.ZN (p_1[15]), .A (slo__sro_n189), .B (n_15));
NOR2_X1 slo__sro_c335 (.ZN (slo__sro_n489), .A1 (p_0[7]), .A2 (Multiplier[7]));
OAI21_X1 slo__sro_c336 (.ZN (slo__sro_n488), .A (slo__sro_n490), .B1 (slo__sro_n491), .B2 (slo__sro_n489));
XNOR2_X1 slo__sro_c337 (.ZN (slo__sro_n487), .A (p_0[7]), .B (Multiplier[7]));
XNOR2_X1 slo__sro_c338 (.ZN (p_1[7]), .A (slo__sro_n487), .B (n_7));
NAND2_X1 slo__sro_c546 (.ZN (slo__sro_n732), .A1 (slo__sro_n190), .A2 (Multiplier[16]));
INV_X1 slo__sro_c174 (.ZN (slo__sro_n251), .A (slo__sro_n488));
NAND2_X1 slo__sro_c175 (.ZN (slo__sro_n250), .A1 (p_0[8]), .A2 (Multiplier[8]));
NOR2_X1 slo__sro_c176 (.ZN (slo__sro_n249), .A1 (p_0[8]), .A2 (Multiplier[8]));
OAI21_X2 slo__sro_c177 (.ZN (slo__sro_n248), .A (slo__sro_n250), .B1 (slo__sro_n251), .B2 (slo__sro_n249));
XNOR2_X1 slo__sro_c178 (.ZN (slo__sro_n247), .A (p_0[8]), .B (Multiplier[8]));
XNOR2_X1 slo__sro_c179 (.ZN (p_1[8]), .A (slo__sro_n247), .B (slo__sro_n488));
INV_X1 slo__xsl_c470 (.ZN (slo__xsl_n643), .A (n_26));
AND2_X2 slo__xsl_c473 (.ZN (n_26), .A1 (CLOCK_slo__sro_n1417), .A2 (slo__sro_n163));
XNOR2_X2 slo__sro_c550 (.ZN (p_1[16]), .A (slo__sro_n729), .B (p_0[16]));
OAI21_X2 slo__sro_c594 (.ZN (slo__sro_n190), .A (slo__sro_n192), .B1 (slo__sro_n193), .B2 (slo__sro_n191));
NOR2_X1 CLOCK_slo__sro_c843 (.ZN (CLOCK_slo__sro_n1108), .A1 (n_1), .A2 (Multiplier[1]));
INV_X1 slo__sro_c312 (.ZN (slo__sro_n468), .A (n_13));
NAND2_X1 slo__sro_c313 (.ZN (slo__sro_n467), .A1 (p_0[13]), .A2 (Multiplier[13]));
NOR2_X1 slo__sro_c314 (.ZN (slo__sro_n466), .A1 (p_0[13]), .A2 (Multiplier[13]));
OAI21_X1 slo__sro_c315 (.ZN (slo__sro_n465), .A (slo__sro_n467), .B1 (slo__sro_n468), .B2 (slo__sro_n466));
XNOR2_X1 slo__sro_c316 (.ZN (slo__sro_n464), .A (p_0[13]), .B (Multiplier[13]));
XNOR2_X1 slo__sro_c317 (.ZN (p_1[13]), .A (n_13), .B (slo__sro_n464));
XNOR2_X1 CLOCK_slo__sro_c845 (.ZN (CLOCK_slo__sro_n1107), .A (n_1), .B (Multiplier[1]));
XNOR2_X1 CLOCK_slo__sro_c846 (.ZN (p_1[1]), .A (CLOCK_slo__sro_n1107), .B (p_0[1]));
NAND2_X1 CLOCK_slo__sro_c869 (.ZN (CLOCK_slo__sro_n1137), .A1 (n_28), .A2 (Multiplier[28]));
NAND2_X1 CLOCK_slo__sro_c870 (.ZN (CLOCK_slo__sro_n1136), .A1 (n_28), .A2 (p_0[28]));
NAND3_X1 CLOCK_slo__sro_c871 (.ZN (n_29), .A1 (CLOCK_slo__sro_n1137), .A2 (CLOCK_slo__sro_n1136), .A3 (CLOCK_slo__sro_n1138));
XNOR2_X1 CLOCK_slo__sro_c872 (.ZN (CLOCK_slo__sro_n1135), .A (p_0[28]), .B (Multiplier[28]));
XNOR2_X1 CLOCK_slo__sro_c873 (.ZN (p_1[28]), .A (CLOCK_slo__sro_n1135), .B (n_28));
NAND2_X1 CLOCK_slo__sro_c919 (.ZN (CLOCK_slo__sro_n1187), .A1 (slo__sro_n248), .A2 (Multiplier[9]));
NAND2_X1 CLOCK_slo__sro_c920 (.ZN (CLOCK_slo__sro_n1186), .A1 (p_0[9]), .A2 (slo__sro_n248));
NAND3_X2 CLOCK_slo__sro_c921 (.ZN (CLOCK_slo__sro_n1185), .A1 (CLOCK_slo__sro_n1186)
    , .A2 (CLOCK_slo__sro_n1187), .A3 (CLOCK_slo__sro_n1188));
XNOR2_X1 CLOCK_slo__sro_c922 (.ZN (CLOCK_slo__sro_n1184), .A (p_0[9]), .B (Multiplier[9]));
XNOR2_X1 CLOCK_slo__sro_c923 (.ZN (p_1[9]), .A (CLOCK_slo__sro_n1184), .B (slo__sro_n248));
NOR2_X1 CLOCK_slo__sro_c1143 (.ZN (CLOCK_slo__sro_n1419), .A1 (p_0[25]), .A2 (Multiplier[25]));
INV_X1 CLOCK_slo__sro_c1144 (.ZN (CLOCK_slo__sro_n1418), .A (CLOCK_slo__sro_n1419));
INV_X1 slo__sro_c648 (.ZN (slo__sro_n864), .A (CLOCK_slo__sro_n1185));
NAND2_X1 slo__sro_c649 (.ZN (slo__sro_n863), .A1 (p_0[10]), .A2 (Multiplier[10]));
NOR2_X1 slo__sro_c650 (.ZN (slo__sro_n862), .A1 (p_0[10]), .A2 (Multiplier[10]));
OAI21_X1 slo__sro_c651 (.ZN (n_11), .A (slo__sro_n863), .B1 (slo__sro_n862), .B2 (slo__sro_n864));
XNOR2_X1 slo__sro_c652 (.ZN (slo__sro_n861), .A (p_0[10]), .B (Multiplier[10]));
XNOR2_X1 slo__sro_c653 (.ZN (p_1[10]), .A (slo__sro_n861), .B (CLOCK_slo__sro_n1185));

endmodule //datapath__0_156

module datapath__0_152 (p_0, p_1, p_2);

output [31:0] p_2;
input [31:0] p_0;
input [31:0] p_1;
wire slo__sro_n808;
wire CLOCK_slo__mro_n1680;
wire n_1;
wire n_2;
wire CLOCK_slo__sro_n1593;
wire n_5;
wire slo__sro_n341;
wire n_7;
wire n_9;
wire n_11;
wire n_13;
wire n_14;
wire n_15;
wire n_16;
wire n_17;
wire slo__sro_n235;
wire n_20;
wire n_21;
wire n_23;
wire n_25;
wire n_26;
wire n_27;
wire n_28;
wire CLOCK_slo__sro_n1592;
wire n_30;
wire n_32;
wire n_0;
wire n_34;
wire n_33;
wire slo__sro_n179;
wire slo__sro_n180;
wire slo__sro_n181;
wire slo__sro_n182;
wire slo__sro_n234;
wire slo__sro_n91;
wire slo__sro_n92;
wire slo__sro_n93;
wire slo__sro_n94;
wire slo__sro_n95;
wire slo__sro_n236;
wire slo__sro_n237;
wire slo__sro_n238;
wire slo__sro_n221;
wire slo__sro_n222;
wire slo__sro_n223;
wire slo__sro_n224;
wire slo__sro_n323;
wire slo__sro_n324;
wire slo__sro_n325;
wire slo__sro_n326;
wire slo__sro_n266;
wire slo__sro_n267;
wire slo__sro_n268;
wire slo__sro_n269;
wire slo__sro_n270;
wire slo__sro_n342;
wire slo__sro_n343;
wire slo__sro_n344;
wire slo__sro_n501;
wire slo__sro_n502;
wire slo__sro_n400;
wire slo__sro_n401;
wire slo__sro_n402;
wire slo__sro_n403;
wire slo__sro_n503;
wire slo__sro_n504;
wire slo__sro_n505;
wire slo__sro_n809;
wire slo__sro_n810;
wire slo__sro_n811;
wire slo__sro_n812;
wire slo__sro_n840;
wire slo__sro_n841;
wire slo__sro_n842;
wire slo__sro_n843;
wire slo__sro_n844;
wire slo__sro_n845;
wire slo__sro_n846;
wire slo__sro_n864;
wire slo__sro_n865;
wire slo__sro_n866;
wire slo__sro_n867;
wire slo__sro_n923;
wire slo__sro_n924;
wire slo__sro_n925;
wire slo__sro_n926;
wire slo__sro_n927;
wire slo__sro_n949;
wire slo__sro_n950;
wire slo__sro_n951;
wire slo__sro_n952;
wire slo__sro_n953;
wire CLOCK_slo__sro_n1548;
wire slo__mro_n985;
wire CLOCK_slo__sro_n1594;
wire CLOCK_slo__sro_n1595;
wire CLOCK_slo__sro_n1633;
wire CLOCK_slo__sro_n1549;
wire CLOCK_slo__sro_n1550;
wire CLOCK_slo__mro_n1561;
wire CLOCK_slo__sro_n1634;
wire CLOCK_slo__sro_n1635;
wire CLOCK_slo__sro_n1636;
wire CLOCK_slo__sro_n1649;
wire CLOCK_slo__sro_n1650;
wire CLOCK_slo__sro_n1651;
wire CLOCK_slo__sro_n1652;
wire CLOCK_slo__sro_n1665;
wire CLOCK_slo__sro_n1666;
wire CLOCK_slo__sro_n1667;
wire CLOCK_slo__sro_n1668;
wire CLOCK_slo__sro_n1669;
wire CLOCK_slo__sro_n1688;
wire CLOCK_slo__sro_n1689;
wire CLOCK_slo__sro_n1690;


INV_X1 i_36 (.ZN (n_34), .A (p_0[30]));
INV_X1 i_35 (.ZN (n_33), .A (p_1[30]));
INV_X1 i_34 (.ZN (n_32), .A (n_30));
XOR2_X1 i_32 (.Z (p_2[31]), .A (p_0[31]), .B (slo__sro_n808));
OAI22_X1 i_31 (.ZN (n_0), .A1 (n_34), .A2 (p_1[30]), .B1 (p_0[30]), .B2 (n_33));
XNOR2_X1 i_0 (.ZN (p_2[30]), .A (n_32), .B (n_0));
INV_X1 slo__sro_c162 (.ZN (slo__sro_n238), .A (p_1[2]));
INV_X1 slo__sro_c667 (.ZN (slo__sro_n867), .A (slo__sro_n235));
FA_X1 i_28 (.CO (n_28), .S (p_2[27]), .A (p_0[27]), .B (p_1[27]), .CI (n_27));
FA_X1 i_27 (.CO (n_27), .S (p_2[26]), .A (p_0[26]), .B (p_1[26]), .CI (n_26));
FA_X1 i_26 (.CO (n_26), .S (p_2[25]), .A (p_0[25]), .B (p_1[25]), .CI (n_25));
FA_X1 i_25 (.CO (n_25), .S (p_2[24]), .A (p_0[24]), .B (p_1[24]), .CI (CLOCK_slo__sro_n1649));
INV_X1 CLOCK_slo__sro_c1264 (.ZN (CLOCK_slo__sro_n1669), .A (n_11));
FA_X1 i_23 (.CO (n_23), .S (p_2[22]), .A (p_0[22]), .B (p_1[22]), .CI (slo__sro_n950));
XNOR2_X2 CLOCK_slo__sro_c1150 (.ZN (CLOCK_slo__sro_n1548), .A (p_1[6]), .B (p_0[6]));
NAND2_X1 slo__sro_c243 (.ZN (slo__sro_n325), .A1 (p_1[9]), .A2 (p_0[9]));
NOR2_X1 slo__sro_c363 (.ZN (slo__sro_n503), .A1 (p_1[18]), .A2 (p_0[18]));
INV_X1 slo__sro_c630 (.ZN (slo__sro_n812), .A (n_30));
NAND2_X1 slo__sro_c163 (.ZN (slo__sro_n237), .A1 (n_2), .A2 (p_0[2]));
FA_X1 i_17 (.CO (n_17), .S (p_2[16]), .A (p_0[16]), .B (p_1[16]), .CI (n_16));
INV_X1 CLOCK_slo__sro_c1236 (.ZN (CLOCK_slo__sro_n1636), .A (n_14));
NAND2_X1 CLOCK_slo__sro_c1250 (.ZN (CLOCK_slo__sro_n1652), .A1 (p_1[23]), .A2 (p_0[23]));
FA_X1 i_14 (.CO (n_14), .S (p_2[13]), .A (p_0[13]), .B (p_1[13]), .CI (n_13));
FA_X1 i_13 (.CO (n_13), .S (p_2[12]), .A (p_0[12]), .B (p_1[12]), .CI (CLOCK_slo__sro_n1666));
XNOR2_X2 CLOCK_slo__mro_c1278 (.ZN (CLOCK_slo__mro_n1680), .A (p_1[23]), .B (p_0[23]));
FA_X1 i_11 (.CO (n_11), .S (p_2[10]), .A (p_0[10]), .B (p_1[10]), .CI (slo__sro_n323));
INV_X1 slo__sro_c258 (.ZN (slo__sro_n344), .A (slo__sro_n502));
BUF_X4 slo__sro_c725 (.Z (slo__sro_n953), .A (n_21));
XNOR2_X2 CLOCK_slo__mro_c1159 (.ZN (CLOCK_slo__mro_n1561), .A (slo__sro_n235), .B (p_0[3]));
NAND2_X1 slo__sro_c259 (.ZN (slo__sro_n343), .A1 (p_1[19]), .A2 (p_0[19]));
FA_X1 i_5 (.CO (n_5), .S (p_2[4]), .A (p_0[4]), .B (p_1[4]), .CI (slo__sro_n864));
INV_X1 slo__sro_c709 (.ZN (slo__sro_n927), .A (n_7));
INV_X1 slo__sro_c242 (.ZN (slo__sro_n326), .A (n_9));
OAI21_X2 slo__sro_c364 (.ZN (slo__sro_n502), .A (slo__sro_n504), .B1 (slo__sro_n505), .B2 (slo__sro_n503));
HA_X1 i_1 (.CO (n_1), .S (p_2[0]), .A (p_0[0]), .B (p_1[0]));
INV_X1 slo__sro_c108 (.ZN (slo__sro_n182), .A (slo__sro_n841));
NAND2_X1 slo__sro_c109 (.ZN (slo__sro_n181), .A1 (p_1[29]), .A2 (p_0[29]));
NOR2_X1 slo__sro_c110 (.ZN (slo__sro_n180), .A1 (p_1[29]), .A2 (p_0[29]));
OAI21_X1 slo__sro_c111 (.ZN (n_30), .A (slo__sro_n181), .B1 (slo__sro_n182), .B2 (slo__sro_n180));
XNOR2_X1 slo__sro_c112 (.ZN (slo__sro_n179), .A (p_1[29]), .B (p_0[29]));
XNOR2_X1 slo__sro_c113 (.ZN (p_2[29]), .A (slo__sro_n841), .B (slo__sro_n179));
INV_X1 slo__sro_c27 (.ZN (slo__sro_n95), .A (n_17));
NAND2_X1 slo__sro_c28 (.ZN (slo__sro_n94), .A1 (p_1[17]), .A2 (p_0[17]));
NOR2_X1 slo__sro_c29 (.ZN (slo__sro_n93), .A1 (p_1[17]), .A2 (p_0[17]));
OAI21_X2 slo__sro_c30 (.ZN (slo__sro_n92), .A (slo__sro_n94), .B1 (slo__sro_n95), .B2 (slo__sro_n93));
XNOR2_X1 slo__sro_c31 (.ZN (slo__sro_n91), .A (p_1[17]), .B (p_0[17]));
XNOR2_X1 slo__sro_c32 (.ZN (p_2[17]), .A (slo__sro_n91), .B (n_17));
NOR2_X2 slo__sro_c164 (.ZN (slo__sro_n236), .A1 (n_2), .A2 (p_0[2]));
OAI21_X2 slo__sro_c165 (.ZN (slo__sro_n235), .A (slo__sro_n237), .B1 (slo__sro_n238), .B2 (slo__sro_n236));
XNOR2_X2 slo__sro_c166 (.ZN (slo__sro_n234), .A (n_2), .B (p_0[2]));
XNOR2_X2 slo__sro_c167 (.ZN (p_2[2]), .A (slo__sro_n234), .B (p_1[2]));
INV_X1 slo__sro_c148 (.ZN (slo__sro_n224), .A (n_20));
NAND2_X1 slo__sro_c149 (.ZN (slo__sro_n223), .A1 (p_1[20]), .A2 (p_0[20]));
NOR2_X1 slo__sro_c150 (.ZN (slo__sro_n222), .A1 (p_1[20]), .A2 (p_0[20]));
OAI21_X1 slo__sro_c151 (.ZN (n_21), .A (slo__sro_n223), .B1 (slo__sro_n224), .B2 (slo__sro_n222));
XNOR2_X1 slo__sro_c152 (.ZN (slo__sro_n221), .A (p_1[20]), .B (p_0[20]));
XNOR2_X1 slo__sro_c153 (.ZN (p_2[20]), .A (slo__sro_n221), .B (n_20));
NOR2_X1 slo__sro_c244 (.ZN (slo__sro_n324), .A1 (p_1[9]), .A2 (p_0[9]));
OAI21_X2 slo__sro_c245 (.ZN (slo__sro_n323), .A (slo__sro_n325), .B1 (slo__sro_n324), .B2 (slo__sro_n326));
NOR2_X1 CLOCK_slo__sro_c1190 (.ZN (CLOCK_slo__sro_n1593), .A1 (p_1[15]), .A2 (p_0[15]));
INV_X1 slo__sro_c189 (.ZN (slo__sro_n270), .A (n_5));
NAND2_X1 slo__sro_c190 (.ZN (slo__sro_n269), .A1 (p_1[5]), .A2 (p_0[5]));
NOR2_X1 slo__sro_c191 (.ZN (slo__sro_n268), .A1 (p_1[5]), .A2 (p_0[5]));
OAI21_X1 slo__sro_c192 (.ZN (slo__sro_n267), .A (slo__sro_n269), .B1 (slo__sro_n270), .B2 (slo__sro_n268));
XNOR2_X2 slo__sro_c193 (.ZN (slo__sro_n266), .A (p_1[5]), .B (p_0[5]));
XNOR2_X2 slo__sro_c194 (.ZN (p_2[5]), .A (slo__sro_n266), .B (n_5));
NOR2_X2 slo__sro_c260 (.ZN (slo__sro_n342), .A1 (p_1[19]), .A2 (p_0[19]));
OAI21_X4 slo__sro_c261 (.ZN (n_20), .A (slo__sro_n343), .B1 (slo__sro_n342), .B2 (slo__sro_n344));
XNOR2_X2 slo__sro_c262 (.ZN (slo__sro_n341), .A (p_1[19]), .B (p_0[19]));
XNOR2_X2 slo__sro_c263 (.ZN (p_2[19]), .A (slo__sro_n341), .B (slo__sro_n502));
INV_X1 slo__sro_c361 (.ZN (slo__sro_n505), .A (slo__sro_n92));
NAND2_X1 slo__sro_c362 (.ZN (slo__sro_n504), .A1 (p_1[18]), .A2 (p_0[18]));
INV_X1 slo__sro_c306 (.ZN (slo__sro_n403), .A (p_1[1]));
NAND2_X1 slo__sro_c307 (.ZN (slo__sro_n402), .A1 (n_1), .A2 (p_0[1]));
NOR2_X1 slo__sro_c308 (.ZN (slo__sro_n401), .A1 (n_1), .A2 (p_0[1]));
OAI21_X2 slo__sro_c309 (.ZN (n_2), .A (slo__sro_n402), .B1 (slo__sro_n403), .B2 (slo__sro_n401));
XNOR2_X2 slo__sro_c310 (.ZN (slo__sro_n400), .A (n_1), .B (p_0[1]));
XNOR2_X1 slo__sro_c311 (.ZN (p_2[1]), .A (slo__sro_n400), .B (p_1[1]));
XNOR2_X2 slo__sro_c365 (.ZN (slo__sro_n501), .A (p_1[18]), .B (p_0[18]));
XNOR2_X2 slo__sro_c366 (.ZN (p_2[18]), .A (slo__sro_n92), .B (slo__sro_n501));
NOR2_X1 slo__sro_c631 (.ZN (slo__sro_n811), .A1 (n_33), .A2 (p_0[30]));
NAND2_X1 slo__sro_c632 (.ZN (slo__sro_n810), .A1 (slo__sro_n811), .A2 (slo__sro_n812));
OR2_X1 slo__sro_c633 (.ZN (slo__sro_n809), .A1 (p_1[30]), .A2 (n_34));
OAI21_X1 slo__sro_c634 (.ZN (slo__sro_n808), .A (slo__sro_n810), .B1 (n_32), .B2 (slo__sro_n809));
INV_X1 slo__sro_c649 (.ZN (slo__sro_n846), .A (p_0[28]));
INV_X1 slo__sro_c650 (.ZN (slo__sro_n845), .A (p_1[28]));
NAND2_X1 slo__sro_c651 (.ZN (slo__sro_n844), .A1 (p_1[28]), .A2 (p_0[28]));
NAND2_X1 slo__sro_c652 (.ZN (slo__sro_n843), .A1 (slo__sro_n845), .A2 (slo__sro_n846));
NAND2_X1 slo__sro_c653 (.ZN (slo__sro_n842), .A1 (n_28), .A2 (slo__sro_n843));
NAND2_X1 slo__sro_c654 (.ZN (slo__sro_n841), .A1 (slo__sro_n842), .A2 (slo__sro_n844));
XNOR2_X1 slo__sro_c655 (.ZN (slo__sro_n840), .A (p_1[28]), .B (p_0[28]));
XNOR2_X1 slo__sro_c656 (.ZN (p_2[28]), .A (n_28), .B (slo__sro_n840));
NAND2_X1 slo__sro_c668 (.ZN (slo__sro_n866), .A1 (p_1[3]), .A2 (p_0[3]));
NOR2_X2 slo__sro_c669 (.ZN (slo__sro_n865), .A1 (p_1[3]), .A2 (p_0[3]));
OAI21_X1 slo__sro_c670 (.ZN (slo__sro_n864), .A (slo__sro_n866), .B1 (slo__sro_n865), .B2 (slo__sro_n867));
INV_X1 CLOCK_slo__sro_c1188 (.ZN (CLOCK_slo__sro_n1595), .A (n_15));
NAND2_X1 CLOCK_slo__sro_c1189 (.ZN (CLOCK_slo__sro_n1594), .A1 (p_1[15]), .A2 (p_0[15]));
NAND2_X1 slo__sro_c710 (.ZN (slo__sro_n926), .A1 (p_1[7]), .A2 (p_0[7]));
NOR2_X1 slo__sro_c711 (.ZN (slo__sro_n925), .A1 (p_1[7]), .A2 (p_0[7]));
OAI21_X1 slo__sro_c712 (.ZN (slo__sro_n924), .A (slo__sro_n926), .B1 (slo__sro_n925), .B2 (slo__sro_n927));
XNOR2_X2 slo__sro_c713 (.ZN (slo__sro_n923), .A (p_1[7]), .B (p_0[7]));
XNOR2_X2 slo__sro_c714 (.ZN (p_2[7]), .A (slo__sro_n923), .B (n_7));
NAND2_X2 slo__sro_c726 (.ZN (slo__sro_n952), .A1 (slo__sro_n953), .A2 (p_0[21]));
OAI21_X4 slo__sro_c727 (.ZN (slo__sro_n951), .A (p_1[21]), .B1 (slo__sro_n953), .B2 (p_0[21]));
NAND2_X2 slo__sro_c728 (.ZN (slo__sro_n950), .A1 (slo__sro_n951), .A2 (slo__sro_n952));
XNOR2_X1 slo__sro_c729 (.ZN (slo__sro_n949), .A (p_1[21]), .B (p_0[21]));
XNOR2_X1 slo__sro_c730 (.ZN (p_2[21]), .A (slo__sro_n949), .B (slo__sro_n953));
XNOR2_X2 CLOCK_slo__sro_c1151 (.ZN (p_2[6]), .A (CLOCK_slo__sro_n1548), .B (slo__sro_n267));
XNOR2_X2 slo__mro_c759 (.ZN (slo__mro_n985), .A (n_9), .B (p_0[9]));
XNOR2_X1 slo__mro_c760 (.ZN (p_2[9]), .A (slo__mro_n985), .B (p_1[9]));
OAI21_X1 CLOCK_slo__sro_c1191 (.ZN (n_16), .A (CLOCK_slo__sro_n1594), .B1 (CLOCK_slo__sro_n1595), .B2 (CLOCK_slo__sro_n1593));
NAND2_X1 CLOCK_slo__sro_c1147 (.ZN (CLOCK_slo__sro_n1550), .A1 (p_1[6]), .A2 (p_0[6]));
OAI21_X1 CLOCK_slo__sro_c1148 (.ZN (CLOCK_slo__sro_n1549), .A (slo__sro_n267), .B1 (p_1[6]), .B2 (p_0[6]));
NAND2_X1 CLOCK_slo__sro_c1149 (.ZN (n_7), .A1 (CLOCK_slo__sro_n1549), .A2 (CLOCK_slo__sro_n1550));
XNOR2_X1 CLOCK_slo__mro_c1160 (.ZN (p_2[3]), .A (CLOCK_slo__mro_n1561), .B (p_1[3]));
XNOR2_X1 CLOCK_slo__sro_c1192 (.ZN (CLOCK_slo__sro_n1592), .A (p_1[15]), .B (p_0[15]));
XNOR2_X1 CLOCK_slo__sro_c1193 (.ZN (p_2[15]), .A (CLOCK_slo__sro_n1592), .B (n_15));
NAND2_X1 CLOCK_slo__sro_c1237 (.ZN (CLOCK_slo__sro_n1635), .A1 (p_1[14]), .A2 (p_0[14]));
NOR2_X1 CLOCK_slo__sro_c1238 (.ZN (CLOCK_slo__sro_n1634), .A1 (p_1[14]), .A2 (p_0[14]));
OAI21_X4 CLOCK_slo__sro_c1239 (.ZN (n_15), .A (CLOCK_slo__sro_n1635), .B1 (CLOCK_slo__sro_n1636), .B2 (CLOCK_slo__sro_n1634));
XNOR2_X1 CLOCK_slo__sro_c1240 (.ZN (CLOCK_slo__sro_n1633), .A (p_1[14]), .B (p_0[14]));
XNOR2_X1 CLOCK_slo__sro_c1241 (.ZN (p_2[14]), .A (CLOCK_slo__sro_n1633), .B (n_14));
NAND2_X1 CLOCK_slo__sro_c1251 (.ZN (CLOCK_slo__sro_n1651), .A1 (n_23), .A2 (p_0[23]));
NAND2_X1 CLOCK_slo__sro_c1252 (.ZN (CLOCK_slo__sro_n1650), .A1 (n_23), .A2 (p_1[23]));
NAND3_X2 CLOCK_slo__sro_c1253 (.ZN (CLOCK_slo__sro_n1649), .A1 (CLOCK_slo__sro_n1651)
    , .A2 (CLOCK_slo__sro_n1650), .A3 (CLOCK_slo__sro_n1652));
NAND2_X1 CLOCK_slo__sro_c1284 (.ZN (CLOCK_slo__sro_n1690), .A1 (slo__sro_n924), .A2 (p_0[8]));
XNOR2_X2 CLOCK_slo__sro_c1255 (.ZN (p_2[23]), .A (CLOCK_slo__mro_n1680), .B (n_23));
NAND2_X1 CLOCK_slo__sro_c1265 (.ZN (CLOCK_slo__sro_n1668), .A1 (p_1[11]), .A2 (p_0[11]));
NOR2_X1 CLOCK_slo__sro_c1266 (.ZN (CLOCK_slo__sro_n1667), .A1 (p_1[11]), .A2 (p_0[11]));
OAI21_X1 CLOCK_slo__sro_c1267 (.ZN (CLOCK_slo__sro_n1666), .A (CLOCK_slo__sro_n1668)
    , .B1 (CLOCK_slo__sro_n1669), .B2 (CLOCK_slo__sro_n1667));
XNOR2_X1 CLOCK_slo__sro_c1268 (.ZN (CLOCK_slo__sro_n1665), .A (p_1[11]), .B (p_0[11]));
XNOR2_X1 CLOCK_slo__sro_c1269 (.ZN (p_2[11]), .A (CLOCK_slo__sro_n1665), .B (n_11));
OAI21_X1 CLOCK_slo__sro_c1285 (.ZN (CLOCK_slo__sro_n1689), .A (p_1[8]), .B1 (slo__sro_n924), .B2 (p_0[8]));
NAND2_X2 CLOCK_slo__sro_c1286 (.ZN (n_9), .A1 (CLOCK_slo__sro_n1689), .A2 (CLOCK_slo__sro_n1690));
XNOR2_X1 CLOCK_slo__sro_c1287 (.ZN (CLOCK_slo__sro_n1688), .A (p_1[8]), .B (p_0[8]));
XNOR2_X1 CLOCK_slo__sro_c1288 (.ZN (p_2[8]), .A (CLOCK_slo__sro_n1688), .B (slo__sro_n924));

endmodule //datapath__0_152

module datapath__0_151 (Multiplier, p_0, p_1);

output [31:0] p_1;
input [31:0] Multiplier;
input [31:0] p_0;
wire CLOCK_slo__mro_n1086;
wire slo__sro_n740;
wire n_1;
wire n_2;
wire n_4;
wire n_5;
wire slo__sro_n785;
wire n_7;
wire n_8;
wire n_9;
wire slo__sro_n446;
wire n_11;
wire n_12;
wire n_13;
wire n_15;
wire n_17;
wire CLOCK_slo__sro_n1134;
wire n_19;
wire n_23;
wire n_27;
wire n_28;
wire n_29;
wire n_30;
wire n_32;
wire n_0;
wire n_34;
wire n_33;
wire n_31;
wire CLOCK_slo__sro_n1131;
wire slo__sro_n72;
wire slo__sro_n73;
wire slo__sro_n74;
wire slo__sro_n75;
wire slo__sro_n88;
wire slo__sro_n89;
wire slo__sro_n90;
wire slo__sro_n91;
wire slo__sro_n92;
wire slo__sro_n120;
wire slo__sro_n121;
wire slo__sro_n122;
wire slo__sro_n123;
wire slo__sro_n137;
wire slo__sro_n138;
wire slo__sro_n139;
wire slo__sro_n140;
wire slo__sro_n154;
wire slo__sro_n155;
wire slo__sro_n156;
wire slo__sro_n157;
wire slo__sro_n158;
wire slo__sro_n171;
wire slo__sro_n172;
wire slo__sro_n173;
wire slo__sro_n174;
wire slo__sro_n175;
wire slo__sro_n191;
wire slo__sro_n192;
wire slo__sro_n193;
wire slo__sro_n194;
wire slo__sro_n209;
wire slo__sro_n210;
wire slo__sro_n211;
wire slo__sro_n212;
wire slo__sro_n248;
wire slo__sro_n249;
wire slo__sro_n250;
wire slo__sro_n251;
wire slo__sro_n252;
wire slo__sro_n490;
wire slo__sro_n444;
wire slo__sro_n445;
wire slo__sro_n280;
wire slo__sro_n281;
wire slo__sro_n282;
wire slo__sro_n283;
wire slo__sro_n284;
wire slo__sro_n447;
wire slo__sro_n491;
wire slo__sro_n492;
wire slo__sro_n493;
wire slo__sro_n494;
wire slo__sro_n741;
wire slo__sro_n742;
wire slo__sro_n743;
wire slo__sro_n744;
wire CLOCK_slo__mro_n1075;
wire CLOCK_slo__sro_n1132;
wire CLOCK_slo__sro_n1133;
wire slo__sro_n782;
wire slo__sro_n783;
wire slo__sro_n784;
wire slo__sro_n594;
wire slo__sro_n595;
wire slo__sro_n596;
wire slo__sro_n597;
wire slo__sro_n598;
wire slo__sro_n786;
wire CLOCK_slo__sro_n1273;
wire CLOCK_slo__sro_n1238;
wire CLOCK_slo__sro_n1239;
wire CLOCK_slo__sro_n1240;
wire CLOCK_slo__sro_n1241;
wire CLOCK_slo__sro_n1274;
wire CLOCK_slo__sro_n1275;
wire CLOCK_slo__sro_n1276;
wire CLOCK_slo__sro_n1277;
wire CLOCK_slo__sro_n1357;
wire CLOCK_slo__sro_n1358;
wire CLOCK_slo__sro_n1359;
wire CLOCK_slo__sro_n1360;


INV_X1 i_36 (.ZN (n_34), .A (Multiplier[30]));
INV_X1 i_35 (.ZN (n_33), .A (p_0[30]));
INV_X1 i_34 (.ZN (n_32), .A (n_30));
OAI33_X1 i_33 (.ZN (n_31), .A1 (n_32), .A2 (p_0[30]), .A3 (n_34), .B1 (n_30), .B2 (n_33), .B3 (Multiplier[30]));
XOR2_X1 i_32 (.Z (p_1[31]), .A (Multiplier[31]), .B (n_31));
OAI22_X1 i_31 (.ZN (n_0), .A1 (n_34), .A2 (p_0[30]), .B1 (Multiplier[30]), .B2 (n_33));
XNOR2_X1 i_0 (.ZN (p_1[30]), .A (n_32), .B (n_0));
INV_X1 slo__sro_c90 (.ZN (slo__sro_n158), .A (n_19));
FA_X1 i_29 (.CO (n_29), .S (p_1[28]), .A (Multiplier[28]), .B (p_0[28]), .CI (n_28));
FA_X1 i_28 (.CO (n_28), .S (p_1[27]), .A (Multiplier[27]), .B (p_0[27]), .CI (n_27));
NAND2_X1 CLOCK_slo__sro_c1046 (.ZN (CLOCK_slo__sro_n1360), .A1 (n_23), .A2 (Multiplier[23]));
INV_X1 slo__sro_c120 (.ZN (slo__sro_n194), .A (n_15));
INV_X1 slo__sro_c55 (.ZN (slo__sro_n123), .A (slo__sro_n191));
FA_X1 i_23 (.CO (n_23), .S (p_1[22]), .A (Multiplier[22]), .B (p_0[22]), .CI (slo__sro_n72));
INV_X1 slo__sro_c28 (.ZN (slo__sro_n92), .A (CLOCK_slo__sro_n1358));
INV_X1 slo__sro_c104 (.ZN (slo__sro_n175), .A (slo__sro_n89));
FA_X1 i_19 (.CO (n_19), .S (p_1[18]), .A (Multiplier[18]), .B (p_0[18]), .CI (slo__sro_n783));
XNOR2_X1 CLOCK_slo__sro_c831 (.ZN (CLOCK_slo__sro_n1131), .A (p_0[6]), .B (Multiplier[6]));
INV_X1 slo__sro_c71 (.ZN (slo__sro_n140), .A (n_29));
INV_X2 slo__sro_c136 (.ZN (slo__sro_n212), .A (slo__sro_n491));
INV_X1 slo__sro_c176 (.ZN (slo__sro_n252), .A (p_0[2]));
NOR2_X1 slo__sro_c564 (.ZN (slo__sro_n742), .A1 (p_0[20]), .A2 (Multiplier[20]));
FA_X1 i_13 (.CO (n_13), .S (p_1[12]), .A (Multiplier[12]), .B (p_0[12]), .CI (n_12));
FA_X1 i_12 (.CO (n_12), .S (p_1[11]), .A (Multiplier[11]), .B (p_0[11]), .CI (n_11));
FA_X1 i_11 (.CO (n_11), .S (p_1[10]), .A (Multiplier[10]), .B (p_0[10]), .CI (slo__sro_n281));
OAI21_X1 slo__sro_c308 (.ZN (n_2), .A (slo__sro_n446), .B1 (slo__sro_n447), .B2 (slo__sro_n445));
NAND2_X1 CLOCK_slo__sro_c977 (.ZN (CLOCK_slo__sro_n1275), .A1 (CLOCK_slo__sro_n1277), .A2 (Multiplier[26]));
FA_X1 i_8 (.CO (n_8), .S (p_1[7]), .A (Multiplier[7]), .B (p_0[7]), .CI (n_7));
BUF_X2 CLOCK_slo__sro_c975 (.Z (CLOCK_slo__sro_n1277), .A (slo__sro_n172));
NAND2_X1 CLOCK_slo__sro_c976 (.ZN (CLOCK_slo__sro_n1276), .A1 (p_0[26]), .A2 (Multiplier[26]));
FA_X1 i_5 (.CO (n_5), .S (p_1[4]), .A (Multiplier[4]), .B (p_0[4]), .CI (n_4));
FA_X1 i_4 (.CO (n_4), .S (p_1[3]), .A (Multiplier[3]), .B (p_0[3]), .CI (slo__sro_n249));
NAND2_X1 slo__sro_c346 (.ZN (slo__sro_n493), .A1 (p_0[13]), .A2 (Multiplier[13]));
NOR2_X1 slo__sro_c347 (.ZN (slo__sro_n492), .A1 (p_0[13]), .A2 (Multiplier[13]));
HA_X1 i_1 (.CO (n_1), .S (p_1[0]), .A (Multiplier[0]), .B (p_0[0]));
INV_X1 slo__sro_c14 (.ZN (slo__sro_n75), .A (slo__sro_n741));
NAND2_X1 slo__sro_c15 (.ZN (slo__sro_n74), .A1 (p_0[21]), .A2 (Multiplier[21]));
NOR2_X1 slo__sro_c16 (.ZN (slo__sro_n73), .A1 (p_0[21]), .A2 (Multiplier[21]));
OAI21_X1 slo__sro_c17 (.ZN (slo__sro_n72), .A (slo__sro_n74), .B1 (slo__sro_n73), .B2 (slo__sro_n75));
INV_X1 CLOCK_slo__sro_c827 (.ZN (CLOCK_slo__sro_n1134), .A (slo__sro_n595));
NAND2_X1 CLOCK_slo__sro_c828 (.ZN (CLOCK_slo__sro_n1133), .A1 (p_0[6]), .A2 (Multiplier[6]));
NAND2_X1 slo__sro_c29 (.ZN (slo__sro_n91), .A1 (p_0[24]), .A2 (Multiplier[24]));
NOR2_X1 slo__sro_c30 (.ZN (slo__sro_n90), .A1 (p_0[24]), .A2 (Multiplier[24]));
OAI21_X1 slo__sro_c31 (.ZN (slo__sro_n89), .A (slo__sro_n91), .B1 (slo__sro_n92), .B2 (slo__sro_n90));
XNOR2_X1 slo__sro_c32 (.ZN (slo__sro_n88), .A (p_0[24]), .B (Multiplier[24]));
XNOR2_X1 slo__sro_c33 (.ZN (p_1[24]), .A (slo__sro_n88), .B (CLOCK_slo__sro_n1358));
NAND2_X1 slo__sro_c56 (.ZN (slo__sro_n122), .A1 (p_0[16]), .A2 (Multiplier[16]));
NOR2_X1 slo__sro_c57 (.ZN (slo__sro_n121), .A1 (p_0[16]), .A2 (Multiplier[16]));
OAI21_X2 slo__sro_c58 (.ZN (n_17), .A (slo__sro_n122), .B1 (slo__sro_n121), .B2 (slo__sro_n123));
XNOR2_X1 slo__sro_c59 (.ZN (slo__sro_n120), .A (p_0[16]), .B (Multiplier[16]));
XNOR2_X1 slo__sro_c60 (.ZN (p_1[16]), .A (slo__sro_n120), .B (slo__sro_n191));
NAND2_X1 slo__sro_c72 (.ZN (slo__sro_n139), .A1 (p_0[29]), .A2 (Multiplier[29]));
NOR2_X1 slo__sro_c73 (.ZN (slo__sro_n138), .A1 (p_0[29]), .A2 (Multiplier[29]));
OAI21_X1 slo__sro_c74 (.ZN (n_30), .A (slo__sro_n139), .B1 (slo__sro_n140), .B2 (slo__sro_n138));
XNOR2_X1 slo__sro_c75 (.ZN (slo__sro_n137), .A (p_0[29]), .B (Multiplier[29]));
XNOR2_X1 slo__sro_c76 (.ZN (p_1[29]), .A (n_29), .B (slo__sro_n137));
NAND2_X1 slo__sro_c91 (.ZN (slo__sro_n157), .A1 (p_0[19]), .A2 (Multiplier[19]));
NOR2_X1 slo__sro_c92 (.ZN (slo__sro_n156), .A1 (p_0[19]), .A2 (Multiplier[19]));
OAI21_X2 slo__sro_c93 (.ZN (slo__sro_n155), .A (slo__sro_n157), .B1 (slo__sro_n158), .B2 (slo__sro_n156));
XNOR2_X1 slo__sro_c94 (.ZN (slo__sro_n154), .A (p_0[19]), .B (Multiplier[19]));
XNOR2_X1 slo__sro_c95 (.ZN (p_1[19]), .A (slo__sro_n154), .B (n_19));
NAND2_X1 slo__sro_c105 (.ZN (slo__sro_n174), .A1 (p_0[25]), .A2 (Multiplier[25]));
NOR2_X2 slo__sro_c106 (.ZN (slo__sro_n173), .A1 (p_0[25]), .A2 (Multiplier[25]));
OAI21_X1 slo__sro_c107 (.ZN (slo__sro_n172), .A (slo__sro_n174), .B1 (slo__sro_n175), .B2 (slo__sro_n173));
XNOR2_X1 slo__sro_c108 (.ZN (slo__sro_n171), .A (p_0[25]), .B (Multiplier[25]));
XNOR2_X1 slo__sro_c109 (.ZN (p_1[25]), .A (slo__sro_n171), .B (slo__sro_n89));
NAND2_X1 slo__sro_c121 (.ZN (slo__sro_n193), .A1 (p_0[15]), .A2 (Multiplier[15]));
NOR2_X1 slo__sro_c122 (.ZN (slo__sro_n192), .A1 (p_0[15]), .A2 (Multiplier[15]));
OAI21_X2 slo__sro_c123 (.ZN (slo__sro_n191), .A (slo__sro_n193), .B1 (slo__sro_n194), .B2 (slo__sro_n192));
XNOR2_X1 CLOCK_slo__mro_c786 (.ZN (CLOCK_slo__mro_n1086), .A (p_0[21]), .B (Multiplier[21]));
XNOR2_X1 CLOCK_slo__mro_c787 (.ZN (p_1[21]), .A (CLOCK_slo__mro_n1086), .B (slo__sro_n741));
NAND2_X1 slo__sro_c137 (.ZN (slo__sro_n211), .A1 (p_0[14]), .A2 (Multiplier[14]));
NOR2_X2 slo__sro_c138 (.ZN (slo__sro_n210), .A1 (p_0[14]), .A2 (Multiplier[14]));
OAI21_X4 slo__sro_c139 (.ZN (n_15), .A (slo__sro_n211), .B1 (slo__sro_n212), .B2 (slo__sro_n210));
XNOR2_X1 slo__sro_c140 (.ZN (slo__sro_n209), .A (p_0[14]), .B (Multiplier[14]));
XNOR2_X1 slo__sro_c141 (.ZN (p_1[14]), .A (slo__sro_n209), .B (slo__sro_n491));
NAND2_X1 slo__sro_c177 (.ZN (slo__sro_n251), .A1 (n_2), .A2 (Multiplier[2]));
NOR2_X1 slo__sro_c178 (.ZN (slo__sro_n250), .A1 (n_2), .A2 (Multiplier[2]));
OAI21_X1 slo__sro_c179 (.ZN (slo__sro_n249), .A (slo__sro_n251), .B1 (slo__sro_n252), .B2 (slo__sro_n250));
XNOR2_X1 slo__sro_c180 (.ZN (slo__sro_n248), .A (n_2), .B (Multiplier[2]));
XNOR2_X1 slo__sro_c181 (.ZN (p_1[2]), .A (slo__sro_n248), .B (p_0[2]));
NAND2_X1 slo__sro_c563 (.ZN (slo__sro_n743), .A1 (p_0[20]), .A2 (Multiplier[20]));
INV_X1 slo__sro_c345 (.ZN (slo__sro_n494), .A (n_13));
INV_X1 slo__sro_c305 (.ZN (slo__sro_n447), .A (p_0[1]));
NAND2_X1 slo__sro_c306 (.ZN (slo__sro_n446), .A1 (n_1), .A2 (Multiplier[1]));
NOR2_X1 slo__sro_c307 (.ZN (slo__sro_n445), .A1 (n_1), .A2 (Multiplier[1]));
INV_X2 slo__sro_c203 (.ZN (slo__sro_n284), .A (n_9));
NAND2_X1 slo__sro_c204 (.ZN (slo__sro_n283), .A1 (p_0[9]), .A2 (Multiplier[9]));
NOR2_X2 slo__sro_c205 (.ZN (slo__sro_n282), .A1 (p_0[9]), .A2 (Multiplier[9]));
OAI21_X2 slo__sro_c206 (.ZN (slo__sro_n281), .A (slo__sro_n283), .B1 (slo__sro_n284), .B2 (slo__sro_n282));
XNOR2_X1 slo__sro_c207 (.ZN (slo__sro_n280), .A (p_0[9]), .B (Multiplier[9]));
XNOR2_X1 slo__sro_c208 (.ZN (p_1[9]), .A (slo__sro_n280), .B (n_9));
XNOR2_X1 slo__sro_c309 (.ZN (slo__sro_n444), .A (n_1), .B (Multiplier[1]));
XNOR2_X1 slo__sro_c310 (.ZN (p_1[1]), .A (p_0[1]), .B (slo__sro_n444));
OAI21_X2 slo__sro_c348 (.ZN (slo__sro_n491), .A (slo__sro_n493), .B1 (slo__sro_n494), .B2 (slo__sro_n492));
XNOR2_X2 slo__sro_c349 (.ZN (slo__sro_n490), .A (p_0[13]), .B (Multiplier[13]));
XNOR2_X2 slo__sro_c350 (.ZN (p_1[13]), .A (slo__sro_n490), .B (n_13));
OAI21_X2 slo__sro_c565 (.ZN (slo__sro_n741), .A (slo__sro_n743), .B1 (slo__sro_n744), .B2 (slo__sro_n742));
XNOR2_X1 slo__sro_c566 (.ZN (slo__sro_n740), .A (p_0[20]), .B (Multiplier[20]));
INV_X1 slo__sro_c562 (.ZN (slo__sro_n744), .A (slo__sro_n155));
XNOR2_X1 slo__sro_c567 (.ZN (p_1[20]), .A (slo__sro_n155), .B (slo__sro_n740));
XNOR2_X2 CLOCK_slo__mro_c778 (.ZN (CLOCK_slo__mro_n1075), .A (n_15), .B (Multiplier[15]));
XNOR2_X2 CLOCK_slo__mro_c779 (.ZN (p_1[15]), .A (CLOCK_slo__mro_n1075), .B (p_0[15]));
NOR2_X1 CLOCK_slo__sro_c829 (.ZN (CLOCK_slo__sro_n1132), .A1 (p_0[6]), .A2 (Multiplier[6]));
OAI21_X1 CLOCK_slo__sro_c830 (.ZN (n_7), .A (CLOCK_slo__sro_n1133), .B1 (CLOCK_slo__sro_n1132), .B2 (CLOCK_slo__sro_n1134));
INV_X1 slo__sro_c597 (.ZN (slo__sro_n786), .A (n_17));
NAND2_X1 slo__sro_c598 (.ZN (slo__sro_n785), .A1 (p_0[17]), .A2 (Multiplier[17]));
NOR2_X2 slo__sro_c599 (.ZN (slo__sro_n784), .A1 (p_0[17]), .A2 (Multiplier[17]));
OAI21_X2 slo__sro_c600 (.ZN (slo__sro_n783), .A (slo__sro_n785), .B1 (slo__sro_n784), .B2 (slo__sro_n786));
XNOR2_X1 slo__sro_c601 (.ZN (slo__sro_n782), .A (p_0[17]), .B (Multiplier[17]));
XNOR2_X1 slo__sro_c602 (.ZN (p_1[17]), .A (slo__sro_n782), .B (n_17));
XNOR2_X1 CLOCK_slo__sro_c832 (.ZN (p_1[6]), .A (CLOCK_slo__sro_n1131), .B (slo__sro_n595));
INV_X1 slo__sro_c438 (.ZN (slo__sro_n598), .A (n_5));
NAND2_X1 slo__sro_c439 (.ZN (slo__sro_n597), .A1 (p_0[5]), .A2 (Multiplier[5]));
NOR2_X1 slo__sro_c440 (.ZN (slo__sro_n596), .A1 (p_0[5]), .A2 (Multiplier[5]));
OAI21_X1 slo__sro_c441 (.ZN (slo__sro_n595), .A (slo__sro_n597), .B1 (slo__sro_n598), .B2 (slo__sro_n596));
XNOR2_X1 slo__sro_c442 (.ZN (slo__sro_n594), .A (p_0[5]), .B (Multiplier[5]));
XNOR2_X1 slo__sro_c443 (.ZN (p_1[5]), .A (slo__sro_n594), .B (n_5));
INV_X1 CLOCK_slo__sro_c942 (.ZN (CLOCK_slo__sro_n1241), .A (n_8));
NAND2_X1 CLOCK_slo__sro_c943 (.ZN (CLOCK_slo__sro_n1240), .A1 (p_0[8]), .A2 (Multiplier[8]));
NOR2_X1 CLOCK_slo__sro_c944 (.ZN (CLOCK_slo__sro_n1239), .A1 (p_0[8]), .A2 (Multiplier[8]));
OAI21_X2 CLOCK_slo__sro_c945 (.ZN (n_9), .A (CLOCK_slo__sro_n1240), .B1 (CLOCK_slo__sro_n1241), .B2 (CLOCK_slo__sro_n1239));
XNOR2_X1 CLOCK_slo__sro_c946 (.ZN (CLOCK_slo__sro_n1238), .A (p_0[8]), .B (Multiplier[8]));
XNOR2_X1 CLOCK_slo__sro_c947 (.ZN (p_1[8]), .A (CLOCK_slo__sro_n1238), .B (n_8));
NAND2_X1 CLOCK_slo__sro_c978 (.ZN (CLOCK_slo__sro_n1274), .A1 (CLOCK_slo__sro_n1277), .A2 (p_0[26]));
NAND3_X2 CLOCK_slo__sro_c979 (.ZN (n_27), .A1 (CLOCK_slo__sro_n1275), .A2 (CLOCK_slo__sro_n1274), .A3 (CLOCK_slo__sro_n1276));
XNOR2_X1 CLOCK_slo__sro_c980 (.ZN (CLOCK_slo__sro_n1273), .A (p_0[26]), .B (Multiplier[26]));
XNOR2_X1 CLOCK_slo__sro_c981 (.ZN (p_1[26]), .A (CLOCK_slo__sro_n1273), .B (CLOCK_slo__sro_n1277));
OAI21_X1 CLOCK_slo__sro_c1047 (.ZN (CLOCK_slo__sro_n1359), .A (p_0[23]), .B1 (n_23), .B2 (Multiplier[23]));
NAND2_X1 CLOCK_slo__sro_c1048 (.ZN (CLOCK_slo__sro_n1358), .A1 (CLOCK_slo__sro_n1359), .A2 (CLOCK_slo__sro_n1360));
XNOR2_X1 CLOCK_slo__sro_c1049 (.ZN (CLOCK_slo__sro_n1357), .A (n_23), .B (Multiplier[23]));
XNOR2_X1 CLOCK_slo__sro_c1050 (.ZN (p_1[23]), .A (CLOCK_slo__sro_n1357), .B (p_0[23]));

endmodule //datapath__0_151

module datapath__0_147 (opt_ipoPP_1, p_0, p_1, p_2);

output [31:0] p_2;
input [31:0] p_0;
input [31:0] p_1;
input opt_ipoPP_1;
wire CLOCK_slo__sro_n1390;
wire n_1;
wire n_2;
wire n_3;
wire n_5;
wire n_6;
wire n_7;
wire n_8;
wire n_9;
wire n_11;
wire n_14;
wire n_15;
wire n_16;
wire n_17;
wire CLOCK_slo__xsl_n1476;
wire slo__sro_n485;
wire n_21;
wire n_22;
wire n_23;
wire n_24;
wire n_25;
wire n_26;
wire n_27;
wire n_29;
wire n_30;
wire n_32;
wire n_0;
wire n_34;
wire n_33;
wire n_31;
wire slo__sro_n118;
wire CLOCK_slo__xsl_n1475;
wire slo__sro_n120;
wire slo__sro_n216;
wire slo__sro_n217;
wire slo__sro_n218;
wire slo__sro_n219;
wire slo__sro_n220;
wire slo__sro_n233;
wire slo__sro_n234;
wire slo__sro_n235;
wire slo__sro_n236;
wire slo__sro_n237;
wire slo__sro_n250;
wire slo__sro_n251;
wire slo__sro_n252;
wire slo__sro_n253;
wire CLOCK_slo__sro_n989;
wire slo__sro_n267;
wire slo__sro_n268;
wire slo__sro_n269;
wire slo__sro_n270;
wire slo__sro_n271;
wire slo__sro_n484;
wire slo__sro_n199;
wire slo__sro_n200;
wire slo__sro_n201;
wire slo__sro_n202;
wire slo__sro_n203;
wire slo__sro_n486;
wire slo__sro_n487;
wire slo__sro_n548;
wire slo__sro_n549;
wire slo__sro_n550;
wire slo__sro_n551;
wire slo__sro_n654;
wire slo__sro_n655;
wire slo__sro_n656;
wire slo__sro_n657;
wire slo__sro_n714;
wire slo__sro_n715;
wire slo__sro_n716;
wire slo__sro_n717;
wire slo__sro_n718;
wire slo__sro_n749;
wire slo__sro_n750;
wire slo__sro_n751;
wire slo__sro_n919;
wire slo__sro_n920;
wire slo__sro_n921;
wire slo__sro_n922;
wire CLOCK_slo__sro_n990;
wire CLOCK_slo__sro_n991;
wire CLOCK_slo__sro_n1016;
wire CLOCK_slo__sro_n1017;
wire CLOCK_slo__sro_n1018;
wire CLOCK_slo__sro_n1019;
wire CLOCK_slo__sro_n1020;
wire CLOCK_slo__sro_n1094;
wire CLOCK_slo__sro_n1095;
wire CLOCK_slo__sro_n1096;
wire CLOCK_slo__sro_n1391;
wire CLOCK_slo__sro_n1303;
wire CLOCK_slo__sro_n1304;
wire CLOCK_slo__sro_n1305;
wire CLOCK_slo__sro_n1306;
wire CLOCK_slo__sro_n1307;


INV_X1 i_36 (.ZN (n_34), .A (p_0[30]));
INV_X1 i_35 (.ZN (n_33), .A (p_1[30]));
INV_X1 i_34 (.ZN (n_32), .A (n_30));
OAI33_X1 i_33 (.ZN (n_31), .A1 (n_32), .A2 (p_1[30]), .A3 (n_34), .B1 (n_30), .B2 (n_33), .B3 (p_0[30]));
XOR2_X1 i_32 (.Z (p_2[31]), .A (p_0[31]), .B (n_31));
OAI22_X1 i_31 (.ZN (n_0), .A1 (n_34), .A2 (p_1[30]), .B1 (p_0[30]), .B2 (n_33));
XNOR2_X1 i_0 (.ZN (p_2[30]), .A (n_32), .B (n_0));
FA_X1 i_30 (.CO (n_30), .S (p_2[29]), .A (p_0[29]), .B (p_1[29]), .CI (n_29));
OR2_X1 CLOCK_slo__sro_c1022 (.ZN (CLOCK_slo__sro_n1391), .A1 (p_1[25]), .A2 (p_0[25]));
NAND2_X1 slo__sro_c529 (.ZN (slo__sro_n751), .A1 (p_1[13]), .A2 (p_0[13]));
FA_X1 i_27 (.CO (n_27), .S (p_2[26]), .A (p_0[26]), .B (p_1[26]), .CI (n_26));
INV_X1 slo__sro_c144 (.ZN (slo__sro_n220), .A (n_9));
FA_X1 i_25 (.CO (n_25), .S (p_2[24]), .A (p_0[24]), .B (p_1[24]), .CI (n_24));
FA_X1 i_24 (.CO (n_24), .S (p_2[23]), .A (p_0[23]), .B (p_1[23]), .CI (n_23));
FA_X1 i_23 (.CO (n_23), .S (p_2[22]), .A (p_0[22]), .B (p_1[22]), .CI (n_22));
NAND2_X1 slo__sro_c451 (.ZN (slo__sro_n657), .A1 (p_1[20]), .A2 (p_0[20]));
INV_X1 slo__sro_c505 (.ZN (slo__sro_n718), .A (n_27));
NAND2_X1 CLOCK_slo__sro_c634 (.ZN (CLOCK_slo__sro_n991), .A1 (p_0[10]), .A2 (p_1[10]));
XNOR2_X1 slo__sro_c342 (.ZN (slo__sro_n484), .A (p_1[14]), .B (p_0[14]));
INV_X1 CLOCK_slo__xsl_c1109 (.ZN (CLOCK_slo__xsl_n1475), .A (CLOCK_slo__xsl_n1476));
FA_X1 i_17 (.CO (n_17), .S (p_2[16]), .A (p_0[16]), .B (p_1[16]), .CI (n_16));
OAI21_X1 CLOCK_slo__sro_c635 (.ZN (CLOCK_slo__sro_n990), .A (slo__sro_n217), .B1 (p_1[10]), .B2 (p_0[10]));
INV_X1 slo__sro_c406 (.ZN (slo__sro_n551), .A (n_21));
INV_X1 slo__sro_c616 (.ZN (slo__sro_n922), .A (p_1[15]));
NAND2_X1 CLOCK_slo__sro_c743 (.ZN (CLOCK_slo__sro_n1096), .A1 (slo__sro_n715), .A2 (p_0[28]));
INV_X1 slo__sro_c338 (.ZN (slo__sro_n487), .A (n_14));
NAND2_X1 CLOCK_slo__sro_c671 (.ZN (CLOCK_slo__sro_n1020), .A1 (p_1[12]), .A2 (p_0[12]));
NAND2_X1 slo__sro_c158 (.ZN (slo__sro_n237), .A1 (p_1[19]), .A2 (p_0[19]));
FA_X1 i_9 (.CO (n_9), .S (p_2[8]), .A (p_0[8]), .B (p_1[8]), .CI (n_8));
FA_X1 i_8 (.CO (n_8), .S (p_2[7]), .A (p_0[7]), .B (p_1[7]), .CI (n_7));
FA_X1 i_7 (.CO (n_7), .S (p_2[6]), .A (p_0[6]), .B (p_1[6]), .CI (n_6));
FA_X1 i_6 (.CO (n_6), .S (p_2[5]), .A (p_0[5]), .B (p_1[5]), .CI (n_5));
FA_X1 i_5 (.CO (n_5), .S (p_2[4]), .A (p_0[4]), .B (p_1[4]), .CI (slo__sro_n251));
INV_X1 slo__sro_c186 (.ZN (slo__sro_n271), .A (n_11));
FA_X1 i_3 (.CO (n_3), .S (p_2[2]), .A (p_0[2]), .B (p_1[2]), .CI (n_2));
FA_X1 i_2 (.CO (n_2), .S (p_2[1]), .A (p_0[1]), .B (p_1[1]), .CI (n_1));
HA_X1 i_1 (.CO (n_1), .S (p_2[0]), .A (p_0[0]), .B (p_1[0]));
NAND2_X1 slo__sro_c53 (.ZN (slo__sro_n120), .A1 (p_0[25]), .A2 (p_1[25]));
INV_X1 CLOCK_slo__xsl_c1108 (.ZN (CLOCK_slo__xsl_n1476), .A (CLOCK_slo__sro_n1304));
NAND2_X1 slo__sro_c55 (.ZN (n_26), .A1 (CLOCK_slo__sro_n1390), .A2 (slo__sro_n120));
XNOR2_X1 slo__sro_c56 (.ZN (slo__sro_n118), .A (p_1[25]), .B (p_0[25]));
XNOR2_X1 slo__sro_c57 (.ZN (p_2[25]), .A (slo__sro_n118), .B (n_25));
NAND2_X1 slo__sro_c145 (.ZN (slo__sro_n219), .A1 (p_1[9]), .A2 (p_0[9]));
NOR2_X1 slo__sro_c146 (.ZN (slo__sro_n218), .A1 (p_1[9]), .A2 (p_0[9]));
OAI21_X2 slo__sro_c147 (.ZN (slo__sro_n217), .A (slo__sro_n219), .B1 (slo__sro_n220), .B2 (slo__sro_n218));
XNOR2_X1 slo__sro_c148 (.ZN (slo__sro_n216), .A (p_1[9]), .B (p_0[9]));
XNOR2_X1 slo__sro_c149 (.ZN (p_2[9]), .A (n_9), .B (slo__sro_n216));
NAND2_X1 slo__sro_c159 (.ZN (slo__sro_n236), .A1 (slo__sro_n200), .A2 (p_0[19]));
NAND2_X1 slo__sro_c160 (.ZN (slo__sro_n235), .A1 (slo__sro_n200), .A2 (p_1[19]));
NAND3_X2 slo__sro_c161 (.ZN (slo__sro_n234), .A1 (slo__sro_n236), .A2 (slo__sro_n235), .A3 (slo__sro_n237));
XNOR2_X1 slo__sro_c162 (.ZN (slo__sro_n233), .A (slo__sro_n200), .B (p_0[19]));
XNOR2_X1 slo__sro_c163 (.ZN (p_2[19]), .A (slo__sro_n233), .B (p_1[19]));
NAND2_X1 slo__sro_c173 (.ZN (slo__sro_n253), .A1 (n_3), .A2 (p_0[3]));
NOR2_X2 slo__sro_c174 (.ZN (slo__sro_n252), .A1 (n_3), .A2 (p_0[3]));
OAI21_X1 slo__sro_c175 (.ZN (slo__sro_n251), .A (slo__sro_n253), .B1 (slo__sro_n252), .B2 (p_1[3]));
XNOR2_X1 slo__sro_c176 (.ZN (slo__sro_n250), .A (n_3), .B (p_0[3]));
XNOR2_X1 slo__sro_c177 (.ZN (p_2[3]), .A (slo__sro_n250), .B (opt_ipoPP_1));
NAND2_X1 slo__sro_c187 (.ZN (slo__sro_n270), .A1 (p_1[11]), .A2 (p_0[11]));
NOR2_X1 slo__sro_c188 (.ZN (slo__sro_n269), .A1 (p_1[11]), .A2 (p_0[11]));
OAI21_X2 slo__sro_c189 (.ZN (slo__sro_n268), .A (slo__sro_n270), .B1 (slo__sro_n271), .B2 (slo__sro_n269));
XNOR2_X2 slo__sro_c190 (.ZN (slo__sro_n267), .A (p_1[11]), .B (p_0[11]));
XNOR2_X2 slo__sro_c191 (.ZN (p_2[11]), .A (slo__sro_n267), .B (n_11));
NAND2_X1 slo__sro_c339 (.ZN (slo__sro_n486), .A1 (p_1[14]), .A2 (p_0[14]));
NOR2_X1 slo__sro_c340 (.ZN (slo__sro_n485), .A1 (p_1[14]), .A2 (p_0[14]));
NAND2_X1 CLOCK_slo__sro_c958 (.ZN (CLOCK_slo__sro_n1306), .A1 (p_1[17]), .A2 (p_0[17]));
INV_X1 slo__sro_c130 (.ZN (slo__sro_n203), .A (CLOCK_slo__sro_n1304));
NAND2_X1 slo__sro_c131 (.ZN (slo__sro_n202), .A1 (p_1[18]), .A2 (p_0[18]));
NOR2_X1 slo__sro_c132 (.ZN (slo__sro_n201), .A1 (p_1[18]), .A2 (p_0[18]));
OAI21_X1 slo__sro_c133 (.ZN (slo__sro_n200), .A (slo__sro_n202), .B1 (slo__sro_n203), .B2 (slo__sro_n201));
XNOR2_X1 slo__sro_c134 (.ZN (slo__sro_n199), .A (p_1[18]), .B (p_0[18]));
XNOR2_X1 slo__sro_c135 (.ZN (p_2[18]), .A (slo__sro_n199), .B (CLOCK_slo__xsl_n1475));
XNOR2_X1 slo__sro_c343 (.ZN (p_2[14]), .A (slo__sro_n484), .B (n_14));
NAND2_X1 slo__sro_c407 (.ZN (slo__sro_n550), .A1 (p_1[21]), .A2 (p_0[21]));
NOR2_X1 slo__sro_c408 (.ZN (slo__sro_n549), .A1 (p_1[21]), .A2 (p_0[21]));
OAI21_X1 slo__sro_c409 (.ZN (n_22), .A (slo__sro_n550), .B1 (slo__sro_n551), .B2 (slo__sro_n549));
XNOR2_X1 slo__sro_c410 (.ZN (slo__sro_n548), .A (p_1[21]), .B (p_0[21]));
XNOR2_X1 slo__sro_c411 (.ZN (p_2[21]), .A (slo__sro_n548), .B (n_21));
NAND2_X1 slo__sro_c452 (.ZN (slo__sro_n656), .A1 (slo__sro_n234), .A2 (p_0[20]));
NAND2_X1 slo__sro_c453 (.ZN (slo__sro_n655), .A1 (slo__sro_n234), .A2 (p_1[20]));
NAND3_X1 slo__sro_c454 (.ZN (n_21), .A1 (slo__sro_n655), .A2 (slo__sro_n657), .A3 (slo__sro_n656));
XNOR2_X1 slo__sro_c455 (.ZN (slo__sro_n654), .A (p_1[20]), .B (p_0[20]));
XNOR2_X1 slo__sro_c456 (.ZN (p_2[20]), .A (slo__sro_n654), .B (slo__sro_n234));
NAND2_X1 slo__sro_c506 (.ZN (slo__sro_n717), .A1 (p_1[27]), .A2 (p_0[27]));
NOR2_X1 slo__sro_c507 (.ZN (slo__sro_n716), .A1 (p_1[27]), .A2 (p_0[27]));
OAI21_X1 slo__sro_c508 (.ZN (slo__sro_n715), .A (slo__sro_n717), .B1 (slo__sro_n718), .B2 (slo__sro_n716));
XNOR2_X1 slo__sro_c509 (.ZN (slo__sro_n714), .A (p_1[27]), .B (p_0[27]));
XNOR2_X1 slo__sro_c510 (.ZN (p_2[27]), .A (n_27), .B (slo__sro_n714));
OAI21_X1 slo__sro_c530 (.ZN (slo__sro_n750), .A (CLOCK_slo__sro_n1017), .B1 (p_1[13]), .B2 (p_0[13]));
NAND2_X1 slo__sro_c531 (.ZN (n_14), .A1 (slo__sro_n750), .A2 (slo__sro_n751));
XNOR2_X2 slo__sro_c532 (.ZN (slo__sro_n749), .A (p_1[13]), .B (p_0[13]));
XNOR2_X1 slo__sro_c533 (.ZN (p_2[13]), .A (slo__sro_n749), .B (CLOCK_slo__sro_n1017));
NAND2_X1 slo__sro_c617 (.ZN (slo__sro_n921), .A1 (n_15), .A2 (p_0[15]));
NOR2_X1 slo__sro_c618 (.ZN (slo__sro_n920), .A1 (n_15), .A2 (p_0[15]));
OAI21_X1 slo__sro_c619 (.ZN (n_16), .A (slo__sro_n921), .B1 (slo__sro_n920), .B2 (slo__sro_n922));
XNOR2_X2 slo__sro_c620 (.ZN (slo__sro_n919), .A (n_15), .B (p_0[15]));
XNOR2_X2 slo__sro_c621 (.ZN (p_2[15]), .A (slo__sro_n919), .B (p_1[15]));
NAND2_X2 CLOCK_slo__sro_c636 (.ZN (n_11), .A1 (CLOCK_slo__sro_n990), .A2 (CLOCK_slo__sro_n991));
XNOR2_X1 CLOCK_slo__sro_c637 (.ZN (CLOCK_slo__sro_n989), .A (slo__sro_n217), .B (p_0[10]));
XNOR2_X1 CLOCK_slo__sro_c638 (.ZN (p_2[10]), .A (CLOCK_slo__sro_n989), .B (p_1[10]));
NAND2_X1 CLOCK_slo__sro_c672 (.ZN (CLOCK_slo__sro_n1019), .A1 (slo__sro_n268), .A2 (p_0[12]));
NAND2_X1 CLOCK_slo__sro_c673 (.ZN (CLOCK_slo__sro_n1018), .A1 (slo__sro_n268), .A2 (p_1[12]));
NAND3_X1 CLOCK_slo__sro_c674 (.ZN (CLOCK_slo__sro_n1017), .A1 (CLOCK_slo__sro_n1020)
    , .A2 (CLOCK_slo__sro_n1018), .A3 (CLOCK_slo__sro_n1019));
XNOR2_X1 CLOCK_slo__sro_c675 (.ZN (CLOCK_slo__sro_n1016), .A (slo__sro_n268), .B (p_0[12]));
XNOR2_X1 CLOCK_slo__sro_c676 (.ZN (p_2[12]), .A (CLOCK_slo__sro_n1016), .B (p_1[12]));
OAI21_X1 CLOCK_slo__sro_c744 (.ZN (CLOCK_slo__sro_n1095), .A (p_1[28]), .B1 (slo__sro_n715), .B2 (p_0[28]));
NAND2_X1 CLOCK_slo__sro_c745 (.ZN (n_29), .A1 (CLOCK_slo__sro_n1095), .A2 (CLOCK_slo__sro_n1096));
XNOR2_X1 CLOCK_slo__sro_c746 (.ZN (CLOCK_slo__sro_n1094), .A (slo__sro_n715), .B (p_0[28]));
XNOR2_X1 CLOCK_slo__sro_c747 (.ZN (p_2[28]), .A (CLOCK_slo__sro_n1094), .B (p_1[28]));
NAND2_X1 CLOCK_slo__sro_c1023 (.ZN (CLOCK_slo__sro_n1390), .A1 (n_25), .A2 (CLOCK_slo__sro_n1391));
INV_X1 CLOCK_slo__sro_c957 (.ZN (CLOCK_slo__sro_n1307), .A (n_17));
OAI21_X2 CLOCK_slo__sro_c880 (.ZN (n_15), .A (slo__sro_n486), .B1 (slo__sro_n485), .B2 (slo__sro_n487));
NOR2_X1 CLOCK_slo__sro_c959 (.ZN (CLOCK_slo__sro_n1305), .A1 (p_1[17]), .A2 (p_0[17]));
OAI21_X1 CLOCK_slo__sro_c960 (.ZN (CLOCK_slo__sro_n1304), .A (CLOCK_slo__sro_n1306)
    , .B1 (CLOCK_slo__sro_n1307), .B2 (CLOCK_slo__sro_n1305));
XNOR2_X1 CLOCK_slo__sro_c961 (.ZN (CLOCK_slo__sro_n1303), .A (p_1[17]), .B (p_0[17]));
XNOR2_X1 CLOCK_slo__sro_c962 (.ZN (p_2[17]), .A (CLOCK_slo__sro_n1303), .B (n_17));

endmodule //datapath__0_147

module datapath__0_146 (opt_ipoPP_1, Multiplier, p_0, p_1);

output [31:0] p_1;
input [31:0] Multiplier;
input [31:0] p_0;
input opt_ipoPP_1;
wire CLOCK_slo__sro_n1258;
wire slo__sro_n472;
wire n_1;
wire n_2;
wire n_3;
wire slo__sro_n374;
wire n_5;
wire n_7;
wire n_8;
wire n_9;
wire n_12;
wire n_13;
wire n_15;
wire n_16;
wire n_17;
wire n_18;
wire n_19;
wire CLOCK_slo__xsl_n1321;
wire n_22;
wire n_23;
wire n_25;
wire n_30;
wire n_32;
wire n_0;
wire n_34;
wire n_33;
wire n_31;
wire slo__sro_n57;
wire slo__sro_n58;
wire slo__sro_n59;
wire slo__sro_n60;
wire slo__sro_n61;
wire slo__sro_n74;
wire slo__sro_n75;
wire slo__sro_n76;
wire slo__sro_n77;
wire slo__sro_n89;
wire slo__sro_n90;
wire slo__sro_n91;
wire slo__sro_n92;
wire slo__sro_n93;
wire slo__sro_n106;
wire slo__sro_n107;
wire slo__sro_n108;
wire slo__sro_n109;
wire slo__sro_n110;
wire slo__sro_n123;
wire slo__sro_n124;
wire slo__sro_n125;
wire slo__sro_n126;
wire slo__sro_n151;
wire slo__sro_n152;
wire slo__sro_n153;
wire slo__sro_n154;
wire slo__sro_n410;
wire slo__sro_n372;
wire slo__sro_n373;
wire slo__sro_n211;
wire slo__sro_n212;
wire slo__sro_n213;
wire slo__sro_n214;
wire CLOCK_slo__mro_n1245;
wire slo__sro_n411;
wire slo__sro_n412;
wire slo__sro_n413;
wire slo__sro_n473;
wire slo__sro_n474;
wire slo__sro_n475;
wire slo__sro_n476;
wire slo__sro_n661;
wire slo__sro_n662;
wire slo__sro_n663;
wire slo__sro_n664;
wire CLOCK_slo__xsl_n1320;
wire slo__sro_n677;
wire slo__sro_n678;
wire slo__sro_n679;
wire slo__sro_n680;
wire slo__sro_n769;
wire slo__sro_n770;
wire slo__sro_n771;
wire slo__sro_n772;
wire slo__sro_n816;
wire slo__sro_n817;
wire slo__sro_n926;
wire slo__sro_n927;
wire slo__sro_n928;
wire slo__sro_n929;
wire slo__sro_n930;
wire slo__sro_n1042;
wire slo__sro_n1043;
wire slo__sro_n1044;
wire slo__sro_n1045;
wire slo__sro_n1046;
wire CLOCK_slo__sro_n1259;
wire CLOCK_slo__sro_n1260;
wire CLOCK_slo__sro_n1261;
wire CLOCK_slo__mro_n1295;
wire CLOCK_slo__mro_n1663;
wire CLOCK_slo__sro_n1359;
wire CLOCK_slo__sro_n1360;
wire CLOCK_slo__sro_n1361;


INV_X1 i_36 (.ZN (n_34), .A (Multiplier[30]));
INV_X1 i_35 (.ZN (n_33), .A (p_0[30]));
INV_X1 i_34 (.ZN (n_32), .A (n_30));
OAI33_X1 i_33 (.ZN (n_31), .A1 (n_32), .A2 (p_0[30]), .A3 (n_34), .B1 (n_30), .B2 (n_33), .B3 (Multiplier[30]));
XOR2_X1 i_32 (.Z (p_1[31]), .A (Multiplier[31]), .B (n_31));
OAI22_X1 i_31 (.ZN (n_0), .A1 (n_34), .A2 (p_0[30]), .B1 (Multiplier[30]), .B2 (n_33));
XNOR2_X1 i_0 (.ZN (p_1[30]), .A (n_32), .B (n_0));
FA_X1 i_30 (.CO (n_30), .S (p_1[29]), .A (Multiplier[29]), .B (p_0[29]), .CI (slo__sro_n677));
NAND2_X1 slo__sro_c561 (.ZN (slo__sro_n772), .A1 (slo__sro_n58), .A2 (Multiplier[27]));
NAND2_X1 slo__sro_c605 (.ZN (slo__sro_n817), .A1 (Multiplier[7]), .A2 (p_0[7]));
INV_X1 slo__sro_c15 (.ZN (slo__sro_n77), .A (n_18));
INV_X2 slo__sro_c45 (.ZN (slo__sro_n110), .A (n_19));
FA_X1 i_25 (.CO (n_25), .S (p_1[24]), .A (Multiplier[24]), .B (p_0[24]), .CI (slo__sro_n927));
INV_X1 slo__sro_c791 (.ZN (slo__sro_n1046), .A (n_13));
NAND2_X1 slo__sro_c86 (.ZN (slo__sro_n154), .A1 (p_0[9]), .A2 (Multiplier[9]));
FA_X1 i_22 (.CO (n_22), .S (p_1[21]), .A (Multiplier[21]), .B (p_0[21]), .CI (slo__sro_n662));
INV_X1 slo__sro_c494 (.ZN (slo__sro_n680), .A (slo__sro_n770));
INV_X1 slo__sro_c59 (.ZN (slo__sro_n126), .A (n_22));
INV_X1 slo__sro_c31 (.ZN (slo__sro_n93), .A (n_25));
NAND2_X1 slo__sro_c326 (.ZN (slo__sro_n475), .A1 (Multiplier[5]), .A2 (p_0[5]));
FA_X1 i_17 (.CO (n_17), .S (p_1[16]), .A (Multiplier[16]), .B (p_0[16]), .CI (n_16));
FA_X1 i_16 (.CO (n_16), .S (p_1[15]), .A (Multiplier[15]), .B (p_0[15]), .CI (n_15));
FA_X1 i_15 (.CO (n_15), .S (p_1[14]), .A (Multiplier[14]), .B (p_0[14]), .CI (slo__sro_n1043));
XNOR2_X1 CLOCK_slo__mro_c903 (.ZN (p_1[9]), .A (CLOCK_slo__mro_n1245), .B (p_0[9]));
FA_X1 i_12 (.CO (n_12), .S (p_1[11]), .A (Multiplier[11]), .B (p_0[11]), .CI (CLOCK_slo__sro_n1259));
XNOR2_X2 CLOCK_slo__mro_c959 (.ZN (CLOCK_slo__mro_n1295), .A (slo__sro_n770), .B (Multiplier[28]));
INV_X1 slo__sro_c325 (.ZN (slo__sro_n476), .A (n_5));
NOR2_X1 slo__sro_c278 (.ZN (slo__sro_n411), .A1 (p_0[17]), .A2 (Multiplier[17]));
XNOR2_X1 slo__mro_c702 (.ZN (p_1[17]), .A (n_17), .B (slo__sro_n410));
FA_X1 i_7 (.CO (n_7), .S (p_1[6]), .A (Multiplier[6]), .B (p_0[6]), .CI (slo__sro_n473));
NAND2_X1 slo__sro_c482 (.ZN (slo__sro_n664), .A1 (p_0[20]), .A2 (Multiplier[20]));
FA_X1 i_5 (.CO (n_5), .S (p_1[4]), .A (Multiplier[4]), .B (p_0[4]), .CI (slo__sro_n212));
XNOR2_X2 slo__sro_c241 (.ZN (slo__sro_n372), .A (p_0[8]), .B (Multiplier[8]));
FA_X1 i_3 (.CO (n_3), .S (p_1[2]), .A (Multiplier[2]), .B (p_0[2]), .CI (n_2));
FA_X1 i_2 (.CO (n_2), .S (p_1[1]), .A (Multiplier[1]), .B (p_0[1]), .CI (n_1));
HA_X1 i_1 (.CO (n_1), .S (p_1[0]), .A (Multiplier[0]), .B (p_0[0]));
INV_X1 slo__sro_c1 (.ZN (slo__sro_n61), .A (slo__sro_n90));
NAND2_X1 slo__sro_c2 (.ZN (slo__sro_n60), .A1 (p_0[26]), .A2 (Multiplier[26]));
NOR2_X2 slo__sro_c3 (.ZN (slo__sro_n59), .A1 (p_0[26]), .A2 (Multiplier[26]));
OAI21_X2 slo__sro_c4 (.ZN (slo__sro_n58), .A (slo__sro_n60), .B1 (slo__sro_n59), .B2 (slo__sro_n61));
XNOR2_X2 slo__sro_c5 (.ZN (slo__sro_n57), .A (p_0[26]), .B (Multiplier[26]));
XNOR2_X2 slo__sro_c6 (.ZN (p_1[26]), .A (slo__sro_n57), .B (CLOCK_slo__xsl_n1320));
NAND2_X1 slo__sro_c16 (.ZN (slo__sro_n76), .A1 (p_0[18]), .A2 (Multiplier[18]));
NOR2_X1 slo__sro_c17 (.ZN (slo__sro_n75), .A1 (p_0[18]), .A2 (Multiplier[18]));
OAI21_X2 slo__sro_c18 (.ZN (n_19), .A (slo__sro_n76), .B1 (slo__sro_n77), .B2 (slo__sro_n75));
XNOR2_X2 slo__sro_c19 (.ZN (slo__sro_n74), .A (p_0[18]), .B (Multiplier[18]));
XNOR2_X2 slo__sro_c20 (.ZN (p_1[18]), .A (slo__sro_n74), .B (n_18));
NAND2_X1 slo__sro_c32 (.ZN (slo__sro_n92), .A1 (p_0[25]), .A2 (Multiplier[25]));
NOR2_X1 slo__sro_c33 (.ZN (slo__sro_n91), .A1 (p_0[25]), .A2 (Multiplier[25]));
OAI21_X1 slo__sro_c34 (.ZN (slo__sro_n90), .A (slo__sro_n92), .B1 (slo__sro_n93), .B2 (slo__sro_n91));
XNOR2_X1 slo__sro_c35 (.ZN (slo__sro_n89), .A (p_0[25]), .B (Multiplier[25]));
XNOR2_X1 slo__sro_c36 (.ZN (p_1[25]), .A (slo__sro_n89), .B (n_25));
NAND2_X1 slo__sro_c46 (.ZN (slo__sro_n109), .A1 (p_0[19]), .A2 (Multiplier[19]));
NOR2_X2 slo__sro_c47 (.ZN (slo__sro_n108), .A1 (p_0[19]), .A2 (Multiplier[19]));
XNOR2_X1 slo__sro_c49 (.ZN (slo__sro_n106), .A (p_0[19]), .B (Multiplier[19]));
XNOR2_X1 slo__sro_c50 (.ZN (p_1[19]), .A (slo__sro_n106), .B (n_19));
NAND2_X1 slo__sro_c60 (.ZN (slo__sro_n125), .A1 (p_0[22]), .A2 (Multiplier[22]));
NOR2_X1 slo__sro_c61 (.ZN (slo__sro_n124), .A1 (p_0[22]), .A2 (Multiplier[22]));
OAI21_X1 slo__sro_c62 (.ZN (n_23), .A (slo__sro_n125), .B1 (slo__sro_n126), .B2 (slo__sro_n124));
XNOR2_X1 slo__sro_c63 (.ZN (slo__sro_n123), .A (p_0[22]), .B (Multiplier[22]));
XNOR2_X1 slo__sro_c64 (.ZN (p_1[22]), .A (n_22), .B (slo__sro_n123));
NAND2_X1 slo__sro_c87 (.ZN (slo__sro_n153), .A1 (n_9), .A2 (Multiplier[9]));
NAND2_X1 slo__sro_c88 (.ZN (slo__sro_n152), .A1 (n_9), .A2 (p_0[9]));
NAND3_X2 slo__sro_c89 (.ZN (slo__sro_n151), .A1 (slo__sro_n154), .A2 (slo__sro_n152), .A3 (slo__sro_n153));
NAND2_X1 CLOCK_slo__sro_c915 (.ZN (CLOCK_slo__sro_n1261), .A1 (p_0[10]), .A2 (Multiplier[10]));
AOI22_X1 CLOCK_slo__sro_c916 (.ZN (CLOCK_slo__sro_n1260), .A1 (p_0[10]), .A2 (slo__sro_n151)
    , .B1 (slo__sro_n151), .B2 (Multiplier[10]));
INV_X1 slo__sro_c276 (.ZN (slo__sro_n413), .A (n_17));
NAND2_X1 slo__sro_c277 (.ZN (slo__sro_n412), .A1 (p_0[17]), .A2 (Multiplier[17]));
XNOR2_X2 CLOCK_slo__mro_c1259 (.ZN (p_1[7]), .A (CLOCK_slo__mro_n1663), .B (n_7));
OAI21_X4 slo__sro_c239 (.ZN (slo__sro_n373), .A (n_8), .B1 (p_0[8]), .B2 (Multiplier[8]));
NAND2_X2 slo__sro_c240 (.ZN (n_9), .A1 (slo__sro_n373), .A2 (slo__sro_n374));
XNOR2_X2 CLOCK_slo__mro_c902 (.ZN (CLOCK_slo__mro_n1245), .A (n_9), .B (Multiplier[9]));
NAND2_X1 slo__sro_c145 (.ZN (slo__sro_n214), .A1 (n_3), .A2 (Multiplier[3]));
NOR2_X1 slo__sro_c146 (.ZN (slo__sro_n213), .A1 (n_3), .A2 (Multiplier[3]));
OAI21_X1 slo__sro_c147 (.ZN (slo__sro_n212), .A (slo__sro_n214), .B1 (p_0[3]), .B2 (slo__sro_n213));
XNOR2_X1 slo__sro_c148 (.ZN (slo__sro_n211), .A (n_3), .B (Multiplier[3]));
XNOR2_X1 slo__sro_c149 (.ZN (p_1[3]), .A (slo__sro_n211), .B (opt_ipoPP_1));
XNOR2_X2 slo__sro_c242 (.ZN (p_1[8]), .A (slo__sro_n372), .B (n_8));
XNOR2_X1 slo__sro_c280 (.ZN (slo__sro_n410), .A (p_0[17]), .B (Multiplier[17]));
INV_X1 slo__sro_c706 (.ZN (slo__sro_n930), .A (n_23));
NOR2_X1 slo__sro_c327 (.ZN (slo__sro_n474), .A1 (p_0[5]), .A2 (Multiplier[5]));
OAI21_X1 slo__sro_c328 (.ZN (slo__sro_n473), .A (slo__sro_n475), .B1 (slo__sro_n474), .B2 (slo__sro_n476));
XNOR2_X1 slo__sro_c329 (.ZN (slo__sro_n472), .A (p_0[5]), .B (Multiplier[5]));
XNOR2_X1 slo__sro_c330 (.ZN (p_1[5]), .A (slo__sro_n472), .B (n_5));
AOI22_X2 slo__sro_c483 (.ZN (slo__sro_n663), .A1 (p_0[20]), .A2 (slo__sro_n107), .B1 (slo__sro_n107), .B2 (Multiplier[20]));
NAND2_X1 slo__sro_c484 (.ZN (slo__sro_n662), .A1 (slo__sro_n663), .A2 (slo__sro_n664));
XNOR2_X2 slo__sro_c485 (.ZN (slo__sro_n661), .A (slo__sro_n107), .B (Multiplier[20]));
XNOR2_X1 slo__sro_c486 (.ZN (p_1[20]), .A (slo__sro_n661), .B (p_0[20]));
NAND2_X1 slo__sro_c495 (.ZN (slo__sro_n679), .A1 (p_0[28]), .A2 (Multiplier[28]));
NOR2_X1 slo__sro_c496 (.ZN (slo__sro_n678), .A1 (p_0[28]), .A2 (Multiplier[28]));
OAI21_X1 slo__sro_c497 (.ZN (slo__sro_n677), .A (slo__sro_n679), .B1 (slo__sro_n678), .B2 (slo__sro_n680));
INV_X1 CLOCK_slo__xsl_c989 (.ZN (CLOCK_slo__xsl_n1321), .A (slo__sro_n90));
INV_X1 CLOCK_slo__xsl_c990 (.ZN (CLOCK_slo__xsl_n1320), .A (CLOCK_slo__xsl_n1321));
OAI21_X2 slo__sro_c562 (.ZN (slo__sro_n771), .A (p_0[27]), .B1 (slo__sro_n58), .B2 (Multiplier[27]));
NAND2_X2 slo__sro_c563 (.ZN (slo__sro_n770), .A1 (slo__sro_n771), .A2 (slo__sro_n772));
XNOR2_X2 slo__sro_c564 (.ZN (slo__sro_n769), .A (slo__sro_n58), .B (Multiplier[27]));
XNOR2_X2 slo__sro_c565 (.ZN (p_1[27]), .A (slo__sro_n769), .B (p_0[27]));
OAI21_X1 slo__sro_c606 (.ZN (slo__sro_n816), .A (n_7), .B1 (p_0[7]), .B2 (Multiplier[7]));
NAND2_X2 slo__sro_c607 (.ZN (n_8), .A1 (slo__sro_n816), .A2 (slo__sro_n817));
NAND2_X1 slo__sro_c707 (.ZN (slo__sro_n929), .A1 (p_0[23]), .A2 (Multiplier[23]));
NOR2_X1 slo__sro_c708 (.ZN (slo__sro_n928), .A1 (p_0[23]), .A2 (Multiplier[23]));
OAI21_X1 slo__sro_c709 (.ZN (slo__sro_n927), .A (slo__sro_n929), .B1 (slo__sro_n930), .B2 (slo__sro_n928));
XNOR2_X2 slo__sro_c710 (.ZN (slo__sro_n926), .A (p_0[23]), .B (Multiplier[23]));
XNOR2_X2 slo__sro_c711 (.ZN (p_1[23]), .A (slo__sro_n926), .B (n_23));
NAND2_X1 slo__sro_c792 (.ZN (slo__sro_n1045), .A1 (p_0[13]), .A2 (Multiplier[13]));
NOR2_X1 slo__sro_c793 (.ZN (slo__sro_n1044), .A1 (p_0[13]), .A2 (Multiplier[13]));
OAI21_X1 slo__sro_c794 (.ZN (slo__sro_n1043), .A (slo__sro_n1045), .B1 (slo__sro_n1044), .B2 (slo__sro_n1046));
XNOR2_X1 slo__sro_c795 (.ZN (slo__sro_n1042), .A (p_0[13]), .B (Multiplier[13]));
XNOR2_X1 slo__sro_c796 (.ZN (p_1[13]), .A (slo__sro_n1042), .B (n_13));
NAND2_X1 CLOCK_slo__sro_c917 (.ZN (CLOCK_slo__sro_n1259), .A1 (CLOCK_slo__sro_n1260), .A2 (CLOCK_slo__sro_n1261));
XNOR2_X2 CLOCK_slo__sro_c918 (.ZN (CLOCK_slo__sro_n1258), .A (slo__sro_n151), .B (Multiplier[10]));
XNOR2_X2 CLOCK_slo__sro_c919 (.ZN (p_1[10]), .A (CLOCK_slo__sro_n1258), .B (p_0[10]));
XNOR2_X1 CLOCK_slo__mro_c960 (.ZN (p_1[28]), .A (CLOCK_slo__mro_n1295), .B (p_0[28]));
NAND2_X1 CLOCK_slo__mro_c940 (.ZN (slo__sro_n374), .A1 (p_0[8]), .A2 (Multiplier[8]));
XNOR2_X2 CLOCK_slo__mro_c1258 (.ZN (CLOCK_slo__mro_n1663), .A (p_0[7]), .B (Multiplier[7]));
NAND2_X1 CLOCK_slo__sro_c1028 (.ZN (CLOCK_slo__sro_n1361), .A1 (p_0[12]), .A2 (Multiplier[12]));
OAI21_X1 CLOCK_slo__sro_c1029 (.ZN (CLOCK_slo__sro_n1360), .A (n_12), .B1 (p_0[12]), .B2 (Multiplier[12]));
NAND2_X2 CLOCK_slo__sro_c1030 (.ZN (n_13), .A1 (CLOCK_slo__sro_n1361), .A2 (CLOCK_slo__sro_n1360));
XNOR2_X1 CLOCK_slo__sro_c1031 (.ZN (CLOCK_slo__sro_n1359), .A (p_0[12]), .B (Multiplier[12]));
XNOR2_X1 CLOCK_slo__sro_c1032 (.ZN (p_1[12]), .A (CLOCK_slo__sro_n1359), .B (n_12));
OAI21_X2 CLOCK_slo__sro_c1207 (.ZN (n_18), .A (slo__sro_n412), .B1 (slo__sro_n413), .B2 (slo__sro_n411));
OAI21_X4 CLOCK_slo__sro_c1179 (.ZN (slo__sro_n107), .A (slo__sro_n109), .B1 (slo__sro_n110), .B2 (slo__sro_n108));

endmodule //datapath__0_146

module datapath__0_142 (p_0, p_1, p_2);

output [31:0] p_2;
input [31:0] p_0;
input [31:0] p_1;
wire slo__sro_n796;
wire CLOCK_slo__sro_n1280;
wire n_1;
wire n_2;
wire n_4;
wire n_5;
wire n_7;
wire n_8;
wire n_9;
wire n_10;
wire n_11;
wire slo__sro_n289;
wire n_13;
wire n_15;
wire n_17;
wire n_18;
wire n_19;
wire n_20;
wire n_21;
wire n_22;
wire n_24;
wire slo__sro_n797;
wire n_26;
wire n_27;
wire n_29;
wire n_30;
wire n_32;
wire n_0;
wire n_34;
wire n_33;
wire slo__sro_n92;
wire slo__sro_n93;
wire slo__sro_n94;
wire slo__sro_n95;
wire slo__sro_n96;
wire slo__sro_n124;
wire slo__sro_n125;
wire slo__sro_n126;
wire slo__sro_n127;
wire CLOCK_slo__sro_n1265;
wire slo__sro_n138;
wire slo__sro_n139;
wire slo__sro_n140;
wire slo__sro_n155;
wire slo__sro_n156;
wire slo__sro_n157;
wire slo__sro_n158;
wire slo__sro_n172;
wire slo__sro_n173;
wire slo__sro_n174;
wire slo__sro_n175;
wire slo__sro_n176;
wire slo__sro_n237;
wire slo__sro_n238;
wire slo__sro_n239;
wire slo__sro_n240;
wire slo__sro_n241;
wire slo__sro_n206;
wire slo__sro_n207;
wire slo__sro_n208;
wire slo__sro_n209;
wire slo__sro_n210;
wire slo__sro_n290;
wire slo__sro_n291;
wire slo__sro_n292;
wire slo__sro_n331;
wire slo__sro_n332;
wire slo__sro_n333;
wire slo__sro_n334;
wire slo__sro_n335;
wire slo__sro_n384;
wire slo__sro_n385;
wire slo__sro_n386;
wire slo__sro_n422;
wire slo__sro_n423;
wire slo__sro_n424;
wire slo__sro_n425;
wire slo__sro_n552;
wire slo__sro_n555;
wire slo__sro_n553;
wire slo__sro_n554;
wire slo__sro_n650;
wire slo__sro_n651;
wire slo__sro_n652;
wire slo__sro_n663;
wire slo__sro_n664;
wire slo__sro_n665;
wire slo__sro_n666;
wire slo__sro_n667;
wire slo__sro_n798;
wire slo__sro_n799;
wire slo__sro_n817;
wire slo__sro_n818;
wire slo__sro_n819;
wire slo__sro_n820;
wire slo__sro_n821;
wire slo__mro_n914;
wire CLOCK_slo__sro_n1266;
wire CLOCK_slo__sro_n1267;
wire CLOCK_slo__sro_n1268;
wire CLOCK_slo__sro_n1269;
wire CLOCK_slo__sro_n1281;
wire CLOCK_slo__sro_n1282;
wire CLOCK_slo__sro_n1283;
wire CLOCK_slo__sro_n1284;
wire CLOCK_slo__sro_n1330;
wire CLOCK_slo__sro_n1331;
wire CLOCK_slo__sro_n1332;
wire CLOCK_slo__sro_n1333;
wire CLOCK_slo__sro_n1334;
wire CLOCK_slo__mro_n1347;
wire CLOCK_slo__sro_n1409;
wire CLOCK_slo__sro_n1410;
wire CLOCK_slo__sro_n1411;
wire CLOCK_slo__sro_n1412;
wire CLOCK_slo__sro_n1474;
wire CLOCK_slo__sro_n1475;
wire CLOCK_slo__sro_n1476;
wire CLOCK_slo__sro_n1477;
wire CLOCK_slo__xsl_n1494;


INV_X1 i_36 (.ZN (n_34), .A (p_0[30]));
INV_X1 i_35 (.ZN (n_33), .A (p_1[30]));
INV_X1 i_34 (.ZN (n_32), .A (n_30));
INV_X1 CLOCK_slo__sro_c857 (.ZN (CLOCK_slo__sro_n1334), .A (n_27));
XOR2_X1 i_32 (.Z (p_2[31]), .A (p_0[31]), .B (CLOCK_slo__sro_n1280));
OAI22_X1 i_31 (.ZN (n_0), .A1 (n_34), .A2 (p_1[30]), .B1 (p_0[30]), .B2 (n_33));
XNOR2_X1 i_0 (.ZN (p_2[30]), .A (n_32), .B (n_0));
FA_X1 i_30 (.CO (n_30), .S (p_2[29]), .A (p_0[29]), .B (p_1[29]), .CI (n_29));
FA_X1 i_29 (.CO (n_29), .S (p_2[28]), .A (p_0[28]), .B (p_1[28]), .CI (CLOCK_slo__sro_n1331));
XNOR2_X1 CLOCK_slo__mro_c871 (.ZN (CLOCK_slo__mro_n1347), .A (p_1[18]), .B (p_0[18]));
FA_X1 i_27 (.CO (n_27), .S (p_2[26]), .A (p_0[26]), .B (p_1[26]), .CI (n_26));
FA_X1 i_26 (.CO (n_26), .S (p_2[25]), .A (p_0[25]), .B (p_1[25]), .CI (slo__sro_n664));
NOR2_X2 slo__sro_c556 (.ZN (slo__sro_n797), .A1 (p_1[6]), .A2 (p_0[6]));
INV_X1 slo__sro_c72 (.ZN (slo__sro_n140), .A (n_8));
INV_X1 slo__sro_c195 (.ZN (slo__sro_n292), .A (p_1[9]));
FA_X1 i_21 (.CO (n_21), .S (p_2[20]), .A (p_0[20]), .B (p_1[20]), .CI (n_20));
FA_X1 i_20 (.CO (n_20), .S (p_2[19]), .A (p_0[19]), .B (p_1[19]), .CI (n_19));
INV_X1 slo__sro_c387 (.ZN (slo__sro_n555), .A (p_1[7]));
FA_X1 i_18 (.CO (n_18), .S (p_2[17]), .A (p_0[17]), .B (p_1[17]), .CI (n_17));
INV_X1 slo__sro_c498 (.ZN (slo__sro_n667), .A (n_24));
INV_X1 slo__sro_c258 (.ZN (slo__sro_n386), .A (n_18));
INV_X1 slo__sro_c105 (.ZN (slo__sro_n176), .A (n_13));
INV_X1 slo__sro_c163 (.ZN (slo__sro_n241), .A (n_22));
XNOR2_X2 slo__mro_c648 (.ZN (slo__mro_n914), .A (n_8), .B (p_0[8]));
NAND2_X1 slo__sro_c196 (.ZN (slo__sro_n291), .A1 (n_9), .A2 (p_0[9]));
NAND2_X1 slo__sro_c388 (.ZN (slo__sro_n554), .A1 (n_7), .A2 (p_0[7]));
NAND2_X1 slo__sro_c225 (.ZN (slo__sro_n334), .A1 (n_15), .A2 (p_0[15]));
INV_X1 slo__sro_c89 (.ZN (slo__sro_n158), .A (slo__sro_n173));
BUF_X2 slo__sro_c575 (.Z (slo__sro_n821), .A (slo__sro_n207));
INV_X1 slo__sro_c58 (.ZN (slo__sro_n127), .A (slo__sro_n238));
FA_X1 i_5 (.CO (n_5), .S (p_2[4]), .A (p_0[4]), .B (p_1[4]), .CI (n_4));
INV_X1 CLOCK_slo__sro_c806 (.ZN (CLOCK_slo__sro_n1284), .A (n_30));
FA_X1 i_2 (.CO (n_2), .S (p_2[1]), .A (p_0[1]), .B (p_1[1]), .CI (n_1));
HA_X1 i_1 (.CO (n_1), .S (p_2[0]), .A (p_0[0]), .B (p_1[0]));
INV_X1 slo__sro_c31 (.ZN (slo__sro_n96), .A (n_5));
NAND2_X1 slo__sro_c32 (.ZN (slo__sro_n95), .A1 (p_1[5]), .A2 (p_0[5]));
NOR2_X1 slo__sro_c33 (.ZN (slo__sro_n94), .A1 (p_1[5]), .A2 (p_0[5]));
OAI21_X1 slo__sro_c34 (.ZN (slo__sro_n93), .A (slo__sro_n95), .B1 (slo__sro_n96), .B2 (slo__sro_n94));
XNOR2_X2 slo__sro_c35 (.ZN (slo__sro_n92), .A (p_1[5]), .B (p_0[5]));
XNOR2_X1 slo__sro_c36 (.ZN (p_2[5]), .A (slo__sro_n92), .B (n_5));
NAND2_X1 slo__sro_c59 (.ZN (slo__sro_n126), .A1 (p_1[23]), .A2 (p_0[23]));
NOR2_X1 slo__sro_c60 (.ZN (slo__sro_n125), .A1 (p_1[23]), .A2 (p_0[23]));
OAI21_X1 slo__sro_c61 (.ZN (n_24), .A (slo__sro_n126), .B1 (slo__sro_n127), .B2 (slo__sro_n125));
XNOR2_X2 slo__sro_c62 (.ZN (slo__sro_n124), .A (p_1[23]), .B (p_0[23]));
XNOR2_X2 slo__sro_c63 (.ZN (p_2[23]), .A (slo__sro_n124), .B (slo__sro_n238));
NAND2_X1 slo__sro_c73 (.ZN (slo__sro_n139), .A1 (p_1[8]), .A2 (p_0[8]));
NOR2_X2 slo__sro_c74 (.ZN (slo__sro_n138), .A1 (p_1[8]), .A2 (p_0[8]));
OAI21_X2 slo__sro_c75 (.ZN (n_9), .A (slo__sro_n139), .B1 (slo__sro_n138), .B2 (slo__sro_n140));
INV_X1 CLOCK_slo__sro_c792 (.ZN (CLOCK_slo__sro_n1269), .A (n_2));
NAND2_X1 CLOCK_slo__sro_c793 (.ZN (CLOCK_slo__sro_n1268), .A1 (p_1[2]), .A2 (p_0[2]));
NAND2_X1 slo__sro_c90 (.ZN (slo__sro_n157), .A1 (p_1[14]), .A2 (p_0[14]));
NOR2_X2 slo__sro_c91 (.ZN (slo__sro_n156), .A1 (p_1[14]), .A2 (p_0[14]));
OAI21_X2 slo__sro_c92 (.ZN (n_15), .A (slo__sro_n157), .B1 (slo__sro_n156), .B2 (slo__sro_n158));
XNOR2_X2 slo__sro_c93 (.ZN (slo__sro_n155), .A (p_1[14]), .B (p_0[14]));
XNOR2_X1 slo__sro_c94 (.ZN (p_2[14]), .A (slo__sro_n155), .B (slo__sro_n173));
NAND2_X1 slo__sro_c106 (.ZN (slo__sro_n175), .A1 (p_1[13]), .A2 (p_0[13]));
NOR2_X1 slo__sro_c107 (.ZN (slo__sro_n174), .A1 (p_1[13]), .A2 (p_0[13]));
OAI21_X2 slo__sro_c108 (.ZN (slo__sro_n173), .A (slo__sro_n175), .B1 (slo__sro_n176), .B2 (slo__sro_n174));
XNOR2_X1 slo__sro_c109 (.ZN (slo__sro_n172), .A (p_1[13]), .B (p_0[13]));
XNOR2_X1 slo__sro_c110 (.ZN (p_2[13]), .A (slo__sro_n172), .B (n_13));
NAND2_X1 slo__sro_c164 (.ZN (slo__sro_n240), .A1 (p_1[22]), .A2 (p_0[22]));
NOR2_X1 slo__sro_c165 (.ZN (slo__sro_n239), .A1 (p_1[22]), .A2 (p_0[22]));
OAI21_X1 slo__sro_c166 (.ZN (slo__sro_n238), .A (slo__sro_n240), .B1 (slo__sro_n241), .B2 (slo__sro_n239));
XNOR2_X1 slo__sro_c167 (.ZN (slo__sro_n237), .A (p_1[22]), .B (p_0[22]));
XNOR2_X1 slo__sro_c168 (.ZN (p_2[22]), .A (n_22), .B (slo__sro_n237));
INV_X1 slo__sro_c134 (.ZN (slo__sro_n210), .A (n_11));
NAND2_X1 slo__sro_c135 (.ZN (slo__sro_n209), .A1 (p_1[11]), .A2 (p_0[11]));
NOR2_X1 slo__sro_c136 (.ZN (slo__sro_n208), .A1 (p_1[11]), .A2 (p_0[11]));
OAI21_X1 slo__sro_c137 (.ZN (slo__sro_n207), .A (slo__sro_n209), .B1 (slo__sro_n208), .B2 (slo__sro_n210));
XNOR2_X1 slo__sro_c138 (.ZN (slo__sro_n206), .A (p_1[11]), .B (p_0[11]));
XNOR2_X1 slo__sro_c139 (.ZN (p_2[11]), .A (slo__sro_n206), .B (n_11));
NOR2_X1 slo__sro_c197 (.ZN (slo__sro_n290), .A1 (n_9), .A2 (p_0[9]));
OAI21_X1 slo__sro_c198 (.ZN (n_10), .A (slo__sro_n291), .B1 (slo__sro_n292), .B2 (slo__sro_n290));
XNOR2_X1 slo__sro_c199 (.ZN (slo__sro_n289), .A (n_9), .B (p_0[9]));
XNOR2_X1 slo__sro_c200 (.ZN (p_2[9]), .A (p_1[9]), .B (slo__sro_n289));
NAND2_X1 slo__sro_c555 (.ZN (slo__sro_n798), .A1 (p_1[6]), .A2 (p_0[6]));
NAND2_X1 slo__sro_c224 (.ZN (slo__sro_n335), .A1 (p_1[15]), .A2 (p_0[15]));
NAND2_X1 slo__sro_c226 (.ZN (slo__sro_n333), .A1 (p_1[15]), .A2 (n_15));
XNOR2_X2 slo__sro_c228 (.ZN (slo__sro_n331), .A (n_15), .B (p_0[15]));
XNOR2_X1 slo__sro_c229 (.ZN (p_2[15]), .A (slo__sro_n331), .B (p_1[15]));
NAND2_X1 slo__sro_c259 (.ZN (slo__sro_n385), .A1 (p_0[18]), .A2 (p_1[18]));
NOR2_X1 slo__sro_c260 (.ZN (slo__sro_n384), .A1 (p_1[18]), .A2 (p_0[18]));
OAI21_X1 slo__sro_c261 (.ZN (n_19), .A (slo__sro_n385), .B1 (slo__sro_n386), .B2 (slo__sro_n384));
INV_X1 CLOCK_slo__sro_c897 (.ZN (CLOCK_slo__sro_n1412), .A (p_1[3]));
INV_X1 slo__sro_c284 (.ZN (slo__sro_n425), .A (p_1[10]));
NAND2_X1 slo__sro_c285 (.ZN (slo__sro_n424), .A1 (n_10), .A2 (p_0[10]));
NOR2_X1 slo__sro_c286 (.ZN (slo__sro_n423), .A1 (n_10), .A2 (p_0[10]));
OAI21_X1 slo__sro_c287 (.ZN (n_11), .A (slo__sro_n424), .B1 (slo__sro_n425), .B2 (slo__sro_n423));
XNOR2_X1 slo__sro_c288 (.ZN (slo__sro_n422), .A (n_10), .B (p_0[10]));
XNOR2_X1 slo__sro_c289 (.ZN (p_2[10]), .A (slo__sro_n422), .B (p_1[10]));
INV_X2 slo__sro_c554 (.ZN (slo__sro_n799), .A (slo__sro_n93));
XNOR2_X2 slo__sro_c392 (.ZN (p_2[7]), .A (p_1[7]), .B (slo__sro_n552));
NOR2_X1 slo__sro_c389 (.ZN (slo__sro_n553), .A1 (n_7), .A2 (p_0[7]));
OAI21_X2 slo__sro_c390 (.ZN (n_8), .A (slo__sro_n554), .B1 (slo__sro_n555), .B2 (slo__sro_n553));
XNOR2_X1 slo__sro_c391 (.ZN (slo__sro_n552), .A (n_7), .B (p_0[7]));
NAND2_X1 slo__sro_c485 (.ZN (slo__sro_n652), .A1 (p_1[16]), .A2 (p_0[16]));
NOR2_X1 slo__sro_c486 (.ZN (slo__sro_n651), .A1 (p_1[16]), .A2 (p_0[16]));
OAI21_X1 slo__sro_c487 (.ZN (n_17), .A (slo__sro_n652), .B1 (slo__sro_n651), .B2 (slo__sro_n332));
XNOR2_X1 slo__sro_c488 (.ZN (slo__sro_n650), .A (p_1[16]), .B (p_0[16]));
XNOR2_X1 slo__sro_c489 (.ZN (p_2[16]), .A (slo__sro_n650), .B (CLOCK_slo__xsl_n1494));
NAND2_X1 slo__sro_c499 (.ZN (slo__sro_n666), .A1 (p_1[24]), .A2 (p_0[24]));
NOR2_X1 slo__sro_c500 (.ZN (slo__sro_n665), .A1 (p_1[24]), .A2 (p_0[24]));
OAI21_X1 slo__sro_c501 (.ZN (slo__sro_n664), .A (slo__sro_n666), .B1 (slo__sro_n667), .B2 (slo__sro_n665));
XNOR2_X1 slo__sro_c502 (.ZN (slo__sro_n663), .A (p_1[24]), .B (p_0[24]));
XNOR2_X1 slo__sro_c503 (.ZN (p_2[24]), .A (slo__sro_n663), .B (n_24));
OAI21_X2 slo__sro_c557 (.ZN (n_7), .A (slo__sro_n798), .B1 (slo__sro_n797), .B2 (slo__sro_n799));
XNOR2_X2 slo__sro_c558 (.ZN (slo__sro_n796), .A (p_1[6]), .B (p_0[6]));
XNOR2_X1 slo__sro_c559 (.ZN (p_2[6]), .A (slo__sro_n796), .B (slo__sro_n93));
NAND2_X1 slo__sro_c576 (.ZN (slo__sro_n820), .A1 (p_1[12]), .A2 (p_0[12]));
NAND2_X1 slo__sro_c577 (.ZN (slo__sro_n819), .A1 (slo__sro_n821), .A2 (p_0[12]));
NAND2_X1 slo__sro_c578 (.ZN (slo__sro_n818), .A1 (slo__sro_n821), .A2 (p_1[12]));
NAND3_X1 slo__sro_c579 (.ZN (n_13), .A1 (slo__sro_n818), .A2 (slo__sro_n819), .A3 (slo__sro_n820));
XNOR2_X2 slo__sro_c580 (.ZN (slo__sro_n817), .A (p_1[12]), .B (p_0[12]));
XNOR2_X2 slo__sro_c581 (.ZN (p_2[12]), .A (slo__sro_n817), .B (slo__sro_n821));
XNOR2_X1 slo__mro_c649 (.ZN (p_2[8]), .A (slo__mro_n914), .B (p_1[8]));
NOR2_X1 CLOCK_slo__sro_c794 (.ZN (CLOCK_slo__sro_n1267), .A1 (p_1[2]), .A2 (p_0[2]));
OAI21_X2 CLOCK_slo__sro_c795 (.ZN (CLOCK_slo__sro_n1266), .A (CLOCK_slo__sro_n1268)
    , .B1 (CLOCK_slo__sro_n1269), .B2 (CLOCK_slo__sro_n1267));
XNOR2_X1 CLOCK_slo__sro_c796 (.ZN (CLOCK_slo__sro_n1265), .A (p_1[2]), .B (p_0[2]));
XNOR2_X2 CLOCK_slo__sro_c797 (.ZN (p_2[2]), .A (CLOCK_slo__sro_n1265), .B (n_2));
NOR2_X1 CLOCK_slo__sro_c807 (.ZN (CLOCK_slo__sro_n1283), .A1 (n_33), .A2 (p_0[30]));
NAND2_X1 CLOCK_slo__sro_c808 (.ZN (CLOCK_slo__sro_n1282), .A1 (CLOCK_slo__sro_n1283), .A2 (CLOCK_slo__sro_n1284));
OR2_X1 CLOCK_slo__sro_c809 (.ZN (CLOCK_slo__sro_n1281), .A1 (p_1[30]), .A2 (n_34));
OAI21_X1 CLOCK_slo__sro_c810 (.ZN (CLOCK_slo__sro_n1280), .A (CLOCK_slo__sro_n1282)
    , .B1 (n_32), .B2 (CLOCK_slo__sro_n1281));
NAND2_X1 CLOCK_slo__sro_c858 (.ZN (CLOCK_slo__sro_n1333), .A1 (p_1[27]), .A2 (p_0[27]));
NOR2_X1 CLOCK_slo__sro_c859 (.ZN (CLOCK_slo__sro_n1332), .A1 (p_1[27]), .A2 (p_0[27]));
OAI21_X1 CLOCK_slo__sro_c860 (.ZN (CLOCK_slo__sro_n1331), .A (CLOCK_slo__sro_n1333)
    , .B1 (CLOCK_slo__sro_n1334), .B2 (CLOCK_slo__sro_n1332));
XNOR2_X1 CLOCK_slo__sro_c861 (.ZN (CLOCK_slo__sro_n1330), .A (p_1[27]), .B (p_0[27]));
XNOR2_X1 CLOCK_slo__sro_c862 (.ZN (p_2[27]), .A (CLOCK_slo__sro_n1330), .B (n_27));
XNOR2_X1 CLOCK_slo__mro_c872 (.ZN (p_2[18]), .A (CLOCK_slo__mro_n1347), .B (n_18));
NAND2_X1 CLOCK_slo__sro_c898 (.ZN (CLOCK_slo__sro_n1411), .A1 (CLOCK_slo__sro_n1266), .A2 (p_0[3]));
NOR2_X1 CLOCK_slo__sro_c899 (.ZN (CLOCK_slo__sro_n1410), .A1 (CLOCK_slo__sro_n1266), .A2 (p_0[3]));
OAI21_X1 CLOCK_slo__sro_c900 (.ZN (n_4), .A (CLOCK_slo__sro_n1411), .B1 (CLOCK_slo__sro_n1410), .B2 (CLOCK_slo__sro_n1412));
XNOR2_X2 CLOCK_slo__sro_c901 (.ZN (CLOCK_slo__sro_n1409), .A (CLOCK_slo__sro_n1266), .B (p_0[3]));
XNOR2_X2 CLOCK_slo__sro_c902 (.ZN (p_2[3]), .A (CLOCK_slo__sro_n1409), .B (p_1[3]));
INV_X1 CLOCK_slo__sro_c945 (.ZN (CLOCK_slo__sro_n1477), .A (n_21));
NAND2_X1 CLOCK_slo__sro_c946 (.ZN (CLOCK_slo__sro_n1476), .A1 (p_1[21]), .A2 (p_0[21]));
NOR2_X1 CLOCK_slo__sro_c947 (.ZN (CLOCK_slo__sro_n1475), .A1 (p_1[21]), .A2 (p_0[21]));
OAI21_X1 CLOCK_slo__sro_c948 (.ZN (n_22), .A (CLOCK_slo__sro_n1476), .B1 (CLOCK_slo__sro_n1477), .B2 (CLOCK_slo__sro_n1475));
XNOR2_X1 CLOCK_slo__sro_c949 (.ZN (CLOCK_slo__sro_n1474), .A (p_1[21]), .B (p_0[21]));
XNOR2_X1 CLOCK_slo__sro_c950 (.ZN (p_2[21]), .A (n_21), .B (CLOCK_slo__sro_n1474));
INV_X1 CLOCK_slo__xsl_c975 (.ZN (CLOCK_slo__xsl_n1494), .A (slo__sro_n332));
AND3_X1 CLOCK_slo__xsl_c978 (.ZN (slo__sro_n332), .A1 (slo__sro_n335), .A2 (slo__sro_n333), .A3 (slo__sro_n334));

endmodule //datapath__0_142

module datapath__0_141 (Multiplier, p_0, p_1);

output [31:0] p_1;
input [31:0] Multiplier;
input [31:0] p_0;
wire CLOCK_slo__sro_n1185;
wire slo__sro_n629;
wire n_1;
wire n_2;
wire n_3;
wire n_4;
wire n_5;
wire n_6;
wire n_7;
wire n_9;
wire n_11;
wire CLOCK_slo__xsl_n1226;
wire n_14;
wire n_15;
wire n_18;
wire n_19;
wire n_20;
wire n_21;
wire n_22;
wire n_23;
wire n_26;
wire n_27;
wire n_28;
wire n_30;
wire n_32;
wire n_0;
wire n_34;
wire n_33;
wire n_31;
wire slo__sro_n59;
wire slo__sro_n60;
wire slo__sro_n61;
wire slo__sro_n62;
wire slo__sro_n72;
wire slo__sro_n73;
wire slo__sro_n74;
wire slo__sro_n75;
wire slo__sro_n172;
wire slo__sro_n173;
wire slo__sro_n174;
wire slo__sro_n175;
wire slo__sro_n176;
wire slo__sro_n221;
wire slo__sro_n222;
wire slo__sro_n223;
wire slo__sro_n224;
wire slo__sro_n225;
wire slo__sro_n361;
wire slo__sro_n362;
wire slo__sro_n363;
wire slo__sro_n364;
wire slo__sro_n405;
wire slo__sro_n406;
wire slo__sro_n407;
wire slo__sro_n408;
wire slo__sro_n470;
wire slo__sro_n471;
wire slo__sro_n472;
wire slo__sro_n473;
wire slo__sro_n474;
wire slo__sro_n630;
wire slo__sro_n631;
wire slo__sro_n632;
wire slo__sro_n633;
wire slo__sro_n715;
wire slo__sro_n716;
wire slo__sro_n717;
wire slo__sro_n718;
wire slo__sro_n719;
wire slo__sro_n740;
wire slo__sro_n741;
wire slo__sro_n742;
wire slo__sro_n743;
wire slo__sro_n744;
wire slo__sro_n822;
wire slo__sro_n823;
wire slo__sro_n824;
wire slo__sro_n833;
wire slo__sro_n834;
wire slo__sro_n835;
wire slo__sro_n836;
wire slo__sro_n837;
wire CLOCK_slo__sro_n1186;
wire CLOCK_slo__sro_n1187;
wire CLOCK_slo__sro_n1188;
wire CLOCK_slo__sro_n1189;
wire CLOCK_slo__xsl_n1227;
wire CLOCK_slo__sro_n1245;
wire CLOCK_slo__sro_n1246;
wire CLOCK_slo__sro_n1247;
wire CLOCK_slo__sro_n1248;
wire CLOCK_slo__mro_n1637;
wire CLOCK_slo__sro_n1607;
wire CLOCK_slo__sro_n1608;
wire CLOCK_slo__sro_n1609;
wire CLOCK_slo__sro_n1447;
wire CLOCK_slo__sro_n1448;
wire CLOCK_slo__sro_n1449;
wire CLOCK_slo__sro_n1450;


INV_X1 i_36 (.ZN (n_34), .A (Multiplier[30]));
INV_X1 i_35 (.ZN (n_33), .A (p_0[30]));
INV_X1 i_34 (.ZN (n_32), .A (n_30));
OAI33_X1 i_33 (.ZN (n_31), .A1 (n_34), .A2 (p_0[30]), .A3 (n_32), .B1 (n_30), .B2 (n_33), .B3 (Multiplier[30]));
XOR2_X1 i_32 (.Z (p_1[31]), .A (Multiplier[31]), .B (n_31));
OAI22_X1 i_31 (.ZN (n_0), .A1 (n_34), .A2 (p_0[30]), .B1 (Multiplier[30]), .B2 (n_33));
XNOR2_X1 i_0 (.ZN (p_1[30]), .A (n_32), .B (n_0));
FA_X1 i_30 (.CO (n_30), .S (p_1[29]), .A (Multiplier[29]), .B (p_0[29]), .CI (slo__sro_n834));
NAND2_X1 CLOCK_slo__sro_c857 (.ZN (CLOCK_slo__sro_n1188), .A1 (p_0[11]), .A2 (Multiplier[11]));
FA_X1 i_28 (.CO (n_28), .S (p_1[27]), .A (Multiplier[27]), .B (p_0[27]), .CI (n_27));
INV_X1 slo__sro_c111 (.ZN (slo__sro_n176), .A (n_23));
FA_X1 i_26 (.CO (n_26), .S (p_1[25]), .A (Multiplier[25]), .B (p_0[25]), .CI (slo__sro_n630));
INV_X1 slo__sro_c520 (.ZN (slo__sro_n719), .A (p_0[16]));
INV_X2 slo__sro_c153 (.ZN (slo__sro_n225), .A (CLOCK_slo__sro_n1186));
INV_X1 slo__sro_c467 (.ZN (slo__sro_n633), .A (slo__sro_n173));
INV_X1 slo__sro_c614 (.ZN (slo__sro_n837), .A (n_28));
INV_X1 slo__sro_c17 (.ZN (slo__sro_n75), .A (n_26));
INV_X1 slo__sro_c335 (.ZN (slo__sro_n474), .A (n_15));
FA_X1 i_18 (.CO (n_18), .S (p_1[17]), .A (Multiplier[17]), .B (p_0[17]), .CI (slo__sro_n716));
INV_X1 slo__sro_c536 (.ZN (slo__sro_n744), .A (n_7));
NAND2_X1 slo__sro_c468 (.ZN (slo__sro_n632), .A1 (p_0[24]), .A2 (Multiplier[24]));
FA_X1 i_15 (.CO (n_15), .S (p_1[14]), .A (Multiplier[14]), .B (p_0[14]), .CI (n_14));
FA_X1 i_14 (.CO (n_14), .S (p_1[13]), .A (Multiplier[13]), .B (p_0[13]), .CI (slo__sro_n222));
NAND2_X1 slo__sro_c336 (.ZN (slo__sro_n473), .A1 (p_0[15]), .A2 (Multiplier[15]));
INV_X1 CLOCK_slo__sro_c909 (.ZN (CLOCK_slo__sro_n1248), .A (p_0[9]));
FA_X1 i_11 (.CO (n_11), .S (p_1[10]), .A (Multiplier[10]), .B (p_0[10]), .CI (CLOCK_slo__sro_n1245));
XNOR2_X1 CLOCK_slo__mro_c1251 (.ZN (CLOCK_slo__mro_n1637), .A (p_0[9]), .B (Multiplier[9]));
FA_X1 i_9 (.CO (n_9), .S (p_1[8]), .A (Multiplier[8]), .B (p_0[8]), .CI (slo__sro_n741));
NAND2_X1 slo__sro_c602 (.ZN (slo__sro_n824), .A1 (n_20), .A2 (Multiplier[20]));
FA_X1 i_7 (.CO (n_7), .S (p_1[6]), .A (Multiplier[6]), .B (p_0[6]), .CI (n_6));
FA_X1 i_5 (.CO (n_5), .S (p_1[4]), .A (Multiplier[4]), .B (p_0[4]), .CI (n_4));
FA_X1 i_4 (.CO (n_4), .S (p_1[3]), .A (Multiplier[3]), .B (p_0[3]), .CI (n_3));
FA_X1 i_3 (.CO (n_3), .S (p_1[2]), .A (Multiplier[2]), .B (p_0[2]), .CI (n_2));
FA_X1 i_2 (.CO (n_2), .S (p_1[1]), .A (Multiplier[1]), .B (p_0[1]), .CI (n_1));
HA_X1 i_1 (.CO (n_1), .S (p_1[0]), .A (Multiplier[0]), .B (p_0[0]));
INV_X2 slo__sro_c3 (.ZN (slo__sro_n62), .A (n_19));
NAND2_X1 slo__sro_c4 (.ZN (slo__sro_n61), .A1 (p_0[19]), .A2 (Multiplier[19]));
NOR2_X1 slo__sro_c5 (.ZN (slo__sro_n60), .A1 (p_0[19]), .A2 (Multiplier[19]));
XNOR2_X1 CLOCK_slo__mro_c1252 (.ZN (p_1[9]), .A (CLOCK_slo__mro_n1637), .B (n_9));
XNOR2_X1 slo__sro_c7 (.ZN (slo__sro_n59), .A (p_0[19]), .B (Multiplier[19]));
XNOR2_X2 slo__sro_c8 (.ZN (p_1[19]), .A (slo__sro_n59), .B (CLOCK_slo__xsl_n1226));
NAND2_X1 slo__sro_c18 (.ZN (slo__sro_n74), .A1 (p_0[26]), .A2 (Multiplier[26]));
NOR2_X1 slo__sro_c19 (.ZN (slo__sro_n73), .A1 (p_0[26]), .A2 (Multiplier[26]));
OAI21_X1 slo__sro_c20 (.ZN (n_27), .A (slo__sro_n74), .B1 (slo__sro_n73), .B2 (slo__sro_n75));
XNOR2_X1 slo__sro_c21 (.ZN (slo__sro_n72), .A (p_0[26]), .B (Multiplier[26]));
XNOR2_X1 slo__sro_c22 (.ZN (p_1[26]), .A (slo__sro_n72), .B (n_26));
NAND2_X1 slo__sro_c112 (.ZN (slo__sro_n175), .A1 (p_0[23]), .A2 (Multiplier[23]));
NOR2_X1 slo__sro_c113 (.ZN (slo__sro_n174), .A1 (p_0[23]), .A2 (Multiplier[23]));
OAI21_X2 slo__sro_c114 (.ZN (slo__sro_n173), .A (slo__sro_n175), .B1 (slo__sro_n174), .B2 (slo__sro_n176));
XNOR2_X2 slo__sro_c115 (.ZN (slo__sro_n172), .A (p_0[23]), .B (Multiplier[23]));
XNOR2_X2 slo__sro_c116 (.ZN (p_1[23]), .A (slo__sro_n172), .B (n_23));
NAND2_X1 slo__sro_c154 (.ZN (slo__sro_n224), .A1 (p_0[12]), .A2 (Multiplier[12]));
NOR2_X1 slo__sro_c155 (.ZN (slo__sro_n223), .A1 (p_0[12]), .A2 (Multiplier[12]));
OAI21_X1 slo__sro_c156 (.ZN (slo__sro_n222), .A (slo__sro_n224), .B1 (slo__sro_n225), .B2 (slo__sro_n223));
XNOR2_X1 slo__sro_c157 (.ZN (slo__sro_n221), .A (p_0[12]), .B (Multiplier[12]));
XNOR2_X1 slo__sro_c158 (.ZN (p_1[12]), .A (CLOCK_slo__sro_n1186), .B (slo__sro_n221));
INV_X1 slo__sro_c261 (.ZN (slo__sro_n364), .A (n_22));
NAND2_X1 slo__sro_c262 (.ZN (slo__sro_n363), .A1 (p_0[22]), .A2 (Multiplier[22]));
NOR2_X1 slo__sro_c263 (.ZN (slo__sro_n362), .A1 (p_0[22]), .A2 (Multiplier[22]));
OAI21_X2 slo__sro_c264 (.ZN (n_23), .A (slo__sro_n363), .B1 (slo__sro_n364), .B2 (slo__sro_n362));
XNOR2_X1 slo__sro_c265 (.ZN (slo__sro_n361), .A (p_0[22]), .B (Multiplier[22]));
XNOR2_X1 slo__sro_c266 (.ZN (p_1[22]), .A (slo__sro_n361), .B (n_22));
INV_X1 slo__sro_c290 (.ZN (slo__sro_n408), .A (n_18));
NAND2_X1 slo__sro_c291 (.ZN (slo__sro_n407), .A1 (p_0[18]), .A2 (Multiplier[18]));
NOR2_X1 slo__sro_c292 (.ZN (slo__sro_n406), .A1 (p_0[18]), .A2 (Multiplier[18]));
OAI21_X2 slo__sro_c293 (.ZN (n_19), .A (slo__sro_n407), .B1 (slo__sro_n408), .B2 (slo__sro_n406));
XNOR2_X1 slo__sro_c294 (.ZN (slo__sro_n405), .A (p_0[18]), .B (Multiplier[18]));
XNOR2_X1 slo__sro_c295 (.ZN (p_1[18]), .A (slo__sro_n405), .B (n_18));
NOR2_X1 slo__sro_c337 (.ZN (slo__sro_n472), .A1 (p_0[15]), .A2 (Multiplier[15]));
OAI21_X2 slo__sro_c338 (.ZN (slo__sro_n471), .A (slo__sro_n473), .B1 (slo__sro_n474), .B2 (slo__sro_n472));
XNOR2_X1 slo__sro_c339 (.ZN (slo__sro_n470), .A (p_0[15]), .B (Multiplier[15]));
XNOR2_X1 slo__sro_c340 (.ZN (p_1[15]), .A (slo__sro_n470), .B (n_15));
NOR2_X1 slo__sro_c469 (.ZN (slo__sro_n631), .A1 (p_0[24]), .A2 (Multiplier[24]));
OAI21_X1 slo__sro_c470 (.ZN (slo__sro_n630), .A (slo__sro_n632), .B1 (slo__sro_n631), .B2 (slo__sro_n633));
XNOR2_X2 slo__sro_c471 (.ZN (slo__sro_n629), .A (p_0[24]), .B (Multiplier[24]));
XNOR2_X2 slo__sro_c472 (.ZN (p_1[24]), .A (slo__sro_n629), .B (slo__sro_n173));
NAND2_X1 slo__sro_c521 (.ZN (slo__sro_n718), .A1 (slo__sro_n471), .A2 (Multiplier[16]));
NOR2_X2 slo__sro_c522 (.ZN (slo__sro_n717), .A1 (slo__sro_n471), .A2 (Multiplier[16]));
OAI21_X2 slo__sro_c523 (.ZN (slo__sro_n716), .A (slo__sro_n718), .B1 (slo__sro_n717), .B2 (slo__sro_n719));
XNOR2_X1 slo__sro_c524 (.ZN (slo__sro_n715), .A (slo__sro_n471), .B (Multiplier[16]));
XNOR2_X1 slo__sro_c525 (.ZN (p_1[16]), .A (slo__sro_n715), .B (p_0[16]));
NAND2_X1 slo__sro_c537 (.ZN (slo__sro_n743), .A1 (p_0[7]), .A2 (Multiplier[7]));
NOR2_X1 slo__sro_c538 (.ZN (slo__sro_n742), .A1 (p_0[7]), .A2 (Multiplier[7]));
OAI21_X1 slo__sro_c539 (.ZN (slo__sro_n741), .A (slo__sro_n743), .B1 (slo__sro_n742), .B2 (slo__sro_n744));
XNOR2_X2 slo__sro_c540 (.ZN (slo__sro_n740), .A (p_0[7]), .B (Multiplier[7]));
XNOR2_X2 slo__sro_c541 (.ZN (p_1[7]), .A (slo__sro_n740), .B (n_7));
OAI21_X1 slo__sro_c603 (.ZN (slo__sro_n823), .A (p_0[20]), .B1 (n_20), .B2 (Multiplier[20]));
NAND2_X1 slo__sro_c604 (.ZN (n_21), .A1 (slo__sro_n823), .A2 (slo__sro_n824));
XNOR2_X2 slo__sro_c605 (.ZN (slo__sro_n822), .A (n_20), .B (Multiplier[20]));
XNOR2_X2 slo__sro_c606 (.ZN (p_1[20]), .A (slo__sro_n822), .B (p_0[20]));
NAND2_X1 slo__sro_c615 (.ZN (slo__sro_n836), .A1 (p_0[28]), .A2 (Multiplier[28]));
NOR2_X1 slo__sro_c616 (.ZN (slo__sro_n835), .A1 (p_0[28]), .A2 (Multiplier[28]));
OAI21_X1 slo__sro_c617 (.ZN (slo__sro_n834), .A (slo__sro_n836), .B1 (slo__sro_n837), .B2 (slo__sro_n835));
XNOR2_X1 slo__sro_c618 (.ZN (slo__sro_n833), .A (p_0[28]), .B (Multiplier[28]));
XNOR2_X1 slo__sro_c619 (.ZN (p_1[28]), .A (slo__sro_n833), .B (n_28));
NOR2_X1 CLOCK_slo__sro_c858 (.ZN (CLOCK_slo__sro_n1187), .A1 (p_0[11]), .A2 (Multiplier[11]));
OAI21_X2 CLOCK_slo__sro_c859 (.ZN (CLOCK_slo__sro_n1186), .A (CLOCK_slo__sro_n1188)
    , .B1 (CLOCK_slo__sro_n1189), .B2 (CLOCK_slo__sro_n1187));
INV_X2 CLOCK_slo__sro_c856 (.ZN (CLOCK_slo__sro_n1189), .A (n_11));
XNOR2_X1 CLOCK_slo__sro_c860 (.ZN (CLOCK_slo__sro_n1185), .A (p_0[11]), .B (Multiplier[11]));
XNOR2_X1 CLOCK_slo__sro_c861 (.ZN (p_1[11]), .A (n_11), .B (CLOCK_slo__sro_n1185));
INV_X1 CLOCK_slo__xsl_c895 (.ZN (CLOCK_slo__xsl_n1227), .A (n_19));
INV_X1 CLOCK_slo__xsl_c896 (.ZN (CLOCK_slo__xsl_n1226), .A (CLOCK_slo__xsl_n1227));
NAND2_X1 CLOCK_slo__sro_c910 (.ZN (CLOCK_slo__sro_n1247), .A1 (n_9), .A2 (Multiplier[9]));
NOR2_X1 CLOCK_slo__sro_c911 (.ZN (CLOCK_slo__sro_n1246), .A1 (n_9), .A2 (Multiplier[9]));
OAI21_X1 CLOCK_slo__sro_c912 (.ZN (CLOCK_slo__sro_n1245), .A (CLOCK_slo__sro_n1247)
    , .B1 (CLOCK_slo__sro_n1246), .B2 (CLOCK_slo__sro_n1248));
NAND2_X1 CLOCK_slo__sro_c1214 (.ZN (CLOCK_slo__sro_n1609), .A1 (p_0[21]), .A2 (Multiplier[21]));
OAI21_X1 CLOCK_slo__sro_c1215 (.ZN (CLOCK_slo__sro_n1608), .A (n_21), .B1 (p_0[21]), .B2 (Multiplier[21]));
OAI21_X2 CLOCK_slo__sro_c1000 (.ZN (n_20), .A (slo__sro_n61), .B1 (slo__sro_n62), .B2 (slo__sro_n60));
NAND2_X1 CLOCK_slo__sro_c1216 (.ZN (n_22), .A1 (CLOCK_slo__sro_n1608), .A2 (CLOCK_slo__sro_n1609));
XNOR2_X1 CLOCK_slo__sro_c1217 (.ZN (CLOCK_slo__sro_n1607), .A (p_0[21]), .B (Multiplier[21]));
XNOR2_X1 CLOCK_slo__sro_c1218 (.ZN (p_1[21]), .A (CLOCK_slo__sro_n1607), .B (n_21));
INV_X1 CLOCK_slo__sro_c1092 (.ZN (CLOCK_slo__sro_n1450), .A (n_5));
NAND2_X1 CLOCK_slo__sro_c1093 (.ZN (CLOCK_slo__sro_n1449), .A1 (p_0[5]), .A2 (Multiplier[5]));
NOR2_X1 CLOCK_slo__sro_c1094 (.ZN (CLOCK_slo__sro_n1448), .A1 (p_0[5]), .A2 (Multiplier[5]));
OAI21_X1 CLOCK_slo__sro_c1095 (.ZN (n_6), .A (CLOCK_slo__sro_n1449), .B1 (CLOCK_slo__sro_n1450), .B2 (CLOCK_slo__sro_n1448));
XNOR2_X1 CLOCK_slo__sro_c1096 (.ZN (CLOCK_slo__sro_n1447), .A (p_0[5]), .B (Multiplier[5]));
XNOR2_X1 CLOCK_slo__sro_c1097 (.ZN (p_1[5]), .A (CLOCK_slo__sro_n1447), .B (n_5));

endmodule //datapath__0_141

module datapath__0_137 (p_0_9_PP_0, p_0, p_1, p_2);

output [31:0] p_2;
input [31:0] p_0;
input [31:0] p_1;
input p_0_9_PP_0;
wire CLOCK_slo__mro_n1421;
wire slo__sro_n556;
wire n_1;
wire n_2;
wire n_3;
wire n_4;
wire n_5;
wire n_6;
wire n_8;
wire n_9;
wire n_11;
wire CLOCK_slo__mro_n1484;
wire n_14;
wire n_16;
wire CLOCK_slo__xsl_n1445;
wire n_18;
wire n_20;
wire n_21;
wire n_23;
wire n_24;
wire n_25;
wire n_27;
wire n_29;
wire n_30;
wire n_32;
wire n_0;
wire n_34;
wire n_33;
wire n_31;
wire slo__sro_n95;
wire slo__sro_n96;
wire slo__sro_n97;
wire slo__sro_n98;
wire slo__sro_n99;
wire slo__sro_n199;
wire slo__sro_n200;
wire slo__sro_n201;
wire slo__sro_n202;
wire slo__sro_n203;
wire slo__sro_n216;
wire slo__sro_n217;
wire slo__sro_n218;
wire slo__sro_n219;
wire slo__sro_n220;
wire slo__sro_n233;
wire slo__sro_n234;
wire slo__sro_n236;
wire slo__sro_n237;
wire slo__sro_n251;
wire slo__sro_n252;
wire slo__sro_n253;
wire slo__sro_n254;
wire slo__sro_n267;
wire slo__sro_n268;
wire slo__sro_n269;
wire slo__sro_n270;
wire slo__sro_n271;
wire slo__sro_n284;
wire slo__sro_n285;
wire slo__sro_n286;
wire slo__sro_n287;
wire slo__sro_n288;
wire CLOCK_slo__xsl_n1444;
wire slo__sro_n302;
wire slo__sro_n303;
wire slo__sro_n304;
wire slo__sro_n316;
wire slo__sro_n317;
wire slo__sro_n318;
wire slo__sro_n319;
wire slo__sro_n320;
wire slo__sro_n333;
wire slo__sro_n334;
wire slo__sro_n335;
wire slo__sro_n336;
wire slo__sro_n337;
wire slo__sro_n352;
wire slo__sro_n353;
wire slo__sro_n354;
wire slo__sro_n355;
wire slo__sro_n500;
wire slo__sro_n501;
wire slo__sro_n502;
wire slo__sro_n503;
wire slo__sro_n537;
wire slo__sro_n538;
wire slo__sro_n539;
wire slo__sro_n540;
wire slo__sro_n557;
wire slo__sro_n558;
wire slo__sro_n559;
wire slo__n651;
wire slo__sro_n922;
wire slo__sro_n923;
wire slo__sro_n924;
wire slo__sro_n925;
wire CLOCK_slo__mro_n1462;
wire CLOCK_slo__sro_n1564;
wire CLOCK_slo__sro_n1565;
wire CLOCK_slo__sro_n1566;
wire CLOCK_slo__sro_n1612;
wire CLOCK_slo__sro_n1613;
wire CLOCK_slo__sro_n1614;
wire CLOCK_slo__sro_n1615;


INV_X1 i_36 (.ZN (n_34), .A (p_0[30]));
INV_X1 i_35 (.ZN (n_33), .A (p_1[30]));
INV_X1 i_34 (.ZN (n_32), .A (n_30));
OAI33_X1 i_33 (.ZN (n_31), .A1 (n_34), .A2 (p_1[30]), .A3 (n_32), .B1 (n_30), .B2 (n_33), .B3 (p_0[30]));
XOR2_X1 i_32 (.Z (p_2[31]), .A (p_0[31]), .B (n_31));
OAI22_X1 i_31 (.ZN (n_0), .A1 (n_34), .A2 (p_1[30]), .B1 (p_0[30]), .B2 (n_33));
XNOR2_X1 i_0 (.ZN (p_2[30]), .A (n_32), .B (n_0));
FA_X1 i_30 (.CO (n_30), .S (p_2[29]), .A (p_0[29]), .B (p_1[29]), .CI (n_29));
OAI21_X1 slo__sro_c376 (.ZN (slo__sro_n558), .A (p_1[18]), .B1 (n_18), .B2 (p_0[18]));
INV_X1 slo__sro_c149 (.ZN (slo__sro_n237), .A (n_11));
FA_X1 i_27 (.CO (n_27), .S (p_2[26]), .A (p_0[26]), .B (p_1[26]), .CI (slo__sro_n96));
INV_X2 slo__sro_c121 (.ZN (slo__sro_n203), .A (n_21));
XNOR2_X1 CLOCK_slo__mro_c883 (.ZN (CLOCK_slo__mro_n1462), .A (slo__sro_n234), .B (p_0[12]));
FA_X1 i_24 (.CO (n_24), .S (p_2[23]), .A (p_0[23]), .B (p_1[23]), .CI (n_23));
FA_X1 i_23 (.CO (n_23), .S (p_2[22]), .A (p_0[22]), .B (p_1[22]), .CI (slo__sro_n200));
INV_X1 slo__sro_c135 (.ZN (slo__sro_n220), .A (n_27));
NAND2_X1 slo__sro_c362 (.ZN (slo__sro_n539), .A1 (p_1[28]), .A2 (p_0[28]));
NAND2_X1 CLOCK_slo__sro_c1014 (.ZN (CLOCK_slo__sro_n1614), .A1 (p_1[3]), .A2 (p_0[3]));
OAI21_X1 CLOCK_slo__mro_c835 (.ZN (slo__n651), .A (slo__sro_n287), .B1 (slo__sro_n288), .B2 (slo__sro_n286));
INV_X1 slo__sro_c219 (.ZN (slo__sro_n320), .A (n_6));
INV_X1 slo__sro_c205 (.ZN (slo__sro_n304), .A (p_1[17]));
FA_X1 i_16 (.CO (n_16), .S (p_2[15]), .A (p_0[15]), .B (p_1[15]), .CI (slo__sro_n334));
INV_X1 slo__sro_c249 (.ZN (slo__sro_n355), .A (p_1[13]));
NAND2_X1 slo__sro_c375 (.ZN (slo__sro_n559), .A1 (n_18), .A2 (p_0[18]));
INV_X1 slo__sro_c177 (.ZN (slo__sro_n271), .A (n_9));
INV_X1 slo__sro_c163 (.ZN (slo__sro_n254), .A (p_1[12]));
FA_X1 i_11 (.CO (n_11), .S (p_2[10]), .A (p_0[10]), .B (p_1[10]), .CI (slo__sro_n268));
INV_X1 slo__sro_c191 (.ZN (slo__sro_n288), .A (n_16));
FA_X1 i_9 (.CO (n_9), .S (p_2[8]), .A (p_0[8]), .B (p_1[8]), .CI (n_8));
FA_X1 i_8 (.CO (n_8), .S (p_2[7]), .A (p_0[7]), .B (p_1[7]), .CI (slo__sro_n317));
INV_X1 slo__sro_c233 (.ZN (slo__sro_n337), .A (n_14));
FA_X1 i_6 (.CO (n_6), .S (p_2[5]), .A (p_0[5]), .B (p_1[5]), .CI (n_5));
FA_X1 i_5 (.CO (n_5), .S (p_2[4]), .A (p_0[4]), .B (p_1[4]), .CI (n_4));
FA_X1 i_3 (.CO (n_3), .S (p_2[2]), .A (p_0[2]), .B (p_1[2]), .CI (n_2));
FA_X1 i_2 (.CO (n_2), .S (p_2[1]), .A (p_0[1]), .B (p_1[1]), .CI (n_1));
HA_X1 i_1 (.CO (n_1), .S (p_2[0]), .A (p_0[0]), .B (p_1[0]));
INV_X1 slo__sro_c29 (.ZN (slo__sro_n99), .A (n_25));
NAND2_X1 slo__sro_c30 (.ZN (slo__sro_n98), .A1 (p_1[25]), .A2 (p_0[25]));
NOR2_X1 slo__sro_c31 (.ZN (slo__sro_n97), .A1 (p_1[25]), .A2 (p_0[25]));
OAI21_X1 slo__sro_c32 (.ZN (slo__sro_n96), .A (slo__sro_n98), .B1 (slo__sro_n99), .B2 (slo__sro_n97));
XNOR2_X2 slo__sro_c33 (.ZN (slo__sro_n95), .A (p_1[25]), .B (p_0[25]));
INV_X1 CLOCK_slo__sro_c1013 (.ZN (CLOCK_slo__sro_n1615), .A (n_3));
NAND2_X1 slo__sro_c122 (.ZN (slo__sro_n202), .A1 (p_1[21]), .A2 (p_0[21]));
NOR2_X2 slo__sro_c123 (.ZN (slo__sro_n201), .A1 (p_1[21]), .A2 (p_0[21]));
OAI21_X2 slo__sro_c124 (.ZN (slo__sro_n200), .A (slo__sro_n202), .B1 (slo__sro_n203), .B2 (slo__sro_n201));
XNOR2_X1 slo__sro_c125 (.ZN (slo__sro_n199), .A (p_1[21]), .B (p_0[21]));
XNOR2_X1 slo__sro_c126 (.ZN (p_2[21]), .A (slo__sro_n199), .B (n_21));
NAND2_X1 slo__sro_c136 (.ZN (slo__sro_n219), .A1 (p_1[27]), .A2 (p_0[27]));
NOR2_X1 slo__sro_c137 (.ZN (slo__sro_n218), .A1 (p_1[27]), .A2 (p_0[27]));
OAI21_X1 slo__sro_c138 (.ZN (slo__sro_n217), .A (slo__sro_n219), .B1 (slo__sro_n218), .B2 (slo__sro_n220));
XNOR2_X1 slo__sro_c139 (.ZN (slo__sro_n216), .A (p_1[27]), .B (p_0[27]));
XNOR2_X1 slo__sro_c140 (.ZN (p_2[27]), .A (slo__sro_n216), .B (n_27));
NAND2_X1 slo__sro_c150 (.ZN (slo__sro_n236), .A1 (p_1[11]), .A2 (p_0[11]));
NAND2_X1 CLOCK_slo__sro_c972 (.ZN (CLOCK_slo__sro_n1566), .A1 (p_1[19]), .A2 (p_0[19]));
OAI21_X2 slo__sro_c152 (.ZN (slo__sro_n234), .A (slo__sro_n236), .B1 (slo__sro_n237), .B2 (CLOCK_slo__mro_n1484));
XNOR2_X1 slo__sro_c153 (.ZN (slo__sro_n233), .A (p_1[11]), .B (p_0[11]));
XNOR2_X1 slo__sro_c154 (.ZN (p_2[11]), .A (slo__sro_n233), .B (n_11));
NAND2_X1 slo__sro_c164 (.ZN (slo__sro_n253), .A1 (slo__sro_n234), .A2 (p_0[12]));
NOR2_X1 slo__sro_c165 (.ZN (slo__sro_n252), .A1 (slo__sro_n234), .A2 (p_0[12]));
OAI21_X1 slo__sro_c166 (.ZN (slo__sro_n251), .A (slo__sro_n253), .B1 (slo__sro_n252), .B2 (slo__sro_n254));
XNOR2_X2 CLOCK_slo__sro_c939 (.ZN (p_2[25]), .A (slo__sro_n95), .B (n_25));
NAND2_X1 slo__sro_c178 (.ZN (slo__sro_n270), .A1 (p_1[9]), .A2 (p_0_9_PP_0));
NOR2_X1 slo__sro_c179 (.ZN (slo__sro_n269), .A1 (p_1[9]), .A2 (p_0[9]));
OAI21_X1 slo__sro_c180 (.ZN (slo__sro_n268), .A (slo__sro_n270), .B1 (slo__sro_n271), .B2 (slo__sro_n269));
XNOR2_X1 slo__sro_c181 (.ZN (slo__sro_n267), .A (p_1[9]), .B (p_0[9]));
XNOR2_X1 slo__sro_c182 (.ZN (p_2[9]), .A (slo__sro_n267), .B (n_9));
NAND2_X1 slo__sro_c192 (.ZN (slo__sro_n287), .A1 (p_1[16]), .A2 (p_0[16]));
NOR2_X1 slo__sro_c193 (.ZN (slo__sro_n286), .A1 (p_1[16]), .A2 (p_0[16]));
OAI21_X1 slo__sro_c194 (.ZN (slo__sro_n285), .A (slo__sro_n287), .B1 (slo__sro_n288), .B2 (slo__sro_n286));
XNOR2_X1 slo__sro_c195 (.ZN (slo__sro_n284), .A (p_1[16]), .B (p_0[16]));
XNOR2_X1 slo__sro_c196 (.ZN (p_2[16]), .A (slo__sro_n284), .B (n_16));
NAND2_X1 slo__sro_c206 (.ZN (slo__sro_n303), .A1 (slo__sro_n285), .A2 (p_0[17]));
NOR2_X1 slo__sro_c207 (.ZN (slo__sro_n302), .A1 (slo__sro_n285), .A2 (p_0[17]));
OAI21_X2 slo__sro_c208 (.ZN (n_18), .A (slo__sro_n303), .B1 (slo__sro_n302), .B2 (slo__sro_n304));
INV_X1 CLOCK_slo__xsl_c865 (.ZN (CLOCK_slo__xsl_n1444), .A (CLOCK_slo__xsl_n1445));
INV_X2 CLOCK_slo__xsl_c864 (.ZN (CLOCK_slo__xsl_n1445), .A (n_14));
NAND2_X1 slo__sro_c220 (.ZN (slo__sro_n319), .A1 (p_1[6]), .A2 (p_0[6]));
NOR2_X1 slo__sro_c221 (.ZN (slo__sro_n318), .A1 (p_1[6]), .A2 (p_0[6]));
OAI21_X1 slo__sro_c222 (.ZN (slo__sro_n317), .A (slo__sro_n319), .B1 (slo__sro_n318), .B2 (slo__sro_n320));
XNOR2_X1 slo__sro_c223 (.ZN (slo__sro_n316), .A (p_1[6]), .B (p_0[6]));
XNOR2_X1 slo__sro_c224 (.ZN (p_2[6]), .A (slo__sro_n316), .B (n_6));
NAND2_X1 slo__sro_c234 (.ZN (slo__sro_n336), .A1 (p_1[14]), .A2 (p_0[14]));
NOR2_X1 slo__sro_c235 (.ZN (slo__sro_n335), .A1 (p_1[14]), .A2 (p_0[14]));
OAI21_X2 slo__sro_c236 (.ZN (slo__sro_n334), .A (slo__sro_n336), .B1 (slo__sro_n337), .B2 (slo__sro_n335));
XNOR2_X2 slo__sro_c237 (.ZN (slo__sro_n333), .A (p_1[14]), .B (p_0[14]));
XNOR2_X2 slo__sro_c238 (.ZN (p_2[14]), .A (slo__sro_n333), .B (CLOCK_slo__xsl_n1444));
NAND2_X1 slo__sro_c250 (.ZN (slo__sro_n354), .A1 (slo__sro_n251), .A2 (p_0[13]));
NOR2_X1 slo__sro_c251 (.ZN (slo__sro_n353), .A1 (slo__sro_n251), .A2 (p_0[13]));
OAI21_X2 slo__sro_c252 (.ZN (n_14), .A (slo__sro_n354), .B1 (slo__sro_n353), .B2 (slo__sro_n355));
XNOR2_X1 slo__sro_c253 (.ZN (slo__sro_n352), .A (slo__sro_n251), .B (p_0[13]));
XNOR2_X1 slo__sro_c254 (.ZN (p_2[13]), .A (slo__sro_n352), .B (p_1[13]));
INV_X1 slo__sro_c361 (.ZN (slo__sro_n540), .A (slo__sro_n217));
INV_X2 slo__sro_c337 (.ZN (slo__sro_n503), .A (n_20));
NAND2_X1 slo__sro_c338 (.ZN (slo__sro_n502), .A1 (p_1[20]), .A2 (p_0[20]));
NOR2_X1 slo__sro_c339 (.ZN (slo__sro_n501), .A1 (p_1[20]), .A2 (p_0[20]));
OAI21_X2 slo__sro_c340 (.ZN (n_21), .A (slo__sro_n502), .B1 (slo__sro_n503), .B2 (slo__sro_n501));
XNOR2_X1 slo__sro_c341 (.ZN (slo__sro_n500), .A (p_1[20]), .B (p_0[20]));
XNOR2_X1 slo__sro_c342 (.ZN (p_2[20]), .A (slo__sro_n500), .B (n_20));
NOR2_X1 slo__sro_c363 (.ZN (slo__sro_n538), .A1 (p_1[28]), .A2 (p_0[28]));
OAI21_X1 slo__sro_c364 (.ZN (n_29), .A (slo__sro_n539), .B1 (slo__sro_n538), .B2 (slo__sro_n540));
XNOR2_X1 slo__sro_c365 (.ZN (slo__sro_n537), .A (p_1[28]), .B (p_0[28]));
XNOR2_X1 slo__sro_c366 (.ZN (p_2[28]), .A (slo__sro_n537), .B (slo__sro_n217));
NAND2_X1 slo__sro_c377 (.ZN (slo__sro_n557), .A1 (slo__sro_n558), .A2 (slo__sro_n559));
XNOR2_X2 slo__sro_c378 (.ZN (slo__sro_n556), .A (n_18), .B (p_0[18]));
XNOR2_X1 slo__sro_c379 (.ZN (p_2[18]), .A (slo__sro_n556), .B (p_1[18]));
INV_X1 slo__sro_c606 (.ZN (slo__sro_n925), .A (n_24));
XNOR2_X1 CLOCK_slo__mro_c836 (.ZN (CLOCK_slo__mro_n1421), .A (slo__n651), .B (p_0[17]));
NAND2_X1 slo__sro_c607 (.ZN (slo__sro_n924), .A1 (p_1[24]), .A2 (p_0[24]));
NOR2_X1 slo__sro_c608 (.ZN (slo__sro_n923), .A1 (p_1[24]), .A2 (p_0[24]));
OAI21_X1 slo__sro_c609 (.ZN (n_25), .A (slo__sro_n924), .B1 (slo__sro_n925), .B2 (slo__sro_n923));
XNOR2_X2 slo__sro_c610 (.ZN (slo__sro_n922), .A (p_1[24]), .B (p_0[24]));
XNOR2_X2 slo__sro_c611 (.ZN (p_2[24]), .A (n_24), .B (slo__sro_n922));
XNOR2_X1 CLOCK_slo__mro_c884 (.ZN (p_2[12]), .A (CLOCK_slo__mro_n1462), .B (p_1[12]));
NOR2_X4 CLOCK_slo__mro_c916 (.ZN (CLOCK_slo__mro_n1484), .A1 (p_1[11]), .A2 (p_0[11]));
XNOR2_X1 slo__sro_c718 (.ZN (p_2[17]), .A (CLOCK_slo__mro_n1421), .B (p_1[17]));
OAI21_X4 CLOCK_slo__sro_c973 (.ZN (CLOCK_slo__sro_n1565), .A (slo__sro_n557), .B1 (p_1[19]), .B2 (p_0[19]));
NAND2_X2 CLOCK_slo__sro_c974 (.ZN (n_20), .A1 (CLOCK_slo__sro_n1565), .A2 (CLOCK_slo__sro_n1566));
XNOR2_X1 CLOCK_slo__sro_c975 (.ZN (CLOCK_slo__sro_n1564), .A (p_1[19]), .B (p_0[19]));
XNOR2_X1 CLOCK_slo__sro_c976 (.ZN (p_2[19]), .A (CLOCK_slo__sro_n1564), .B (slo__sro_n557));
NOR2_X1 CLOCK_slo__sro_c1015 (.ZN (CLOCK_slo__sro_n1613), .A1 (p_1[3]), .A2 (p_0[3]));
OAI21_X2 CLOCK_slo__sro_c1016 (.ZN (n_4), .A (CLOCK_slo__sro_n1614), .B1 (CLOCK_slo__sro_n1615), .B2 (CLOCK_slo__sro_n1613));
XNOR2_X2 CLOCK_slo__sro_c1017 (.ZN (CLOCK_slo__sro_n1612), .A (p_1[3]), .B (p_0[3]));
XNOR2_X2 CLOCK_slo__sro_c1018 (.ZN (p_2[3]), .A (CLOCK_slo__sro_n1612), .B (n_3));

endmodule //datapath__0_137

module datapath__0_136 (Multiplier, p_0, p_1);

output [31:0] p_1;
input [31:0] Multiplier;
input [31:0] p_0;
wire CLOCK_slo__sro_n1252;
wire slo__sro_n322;
wire n_1;
wire n_2;
wire n_3;
wire n_4;
wire n_5;
wire n_6;
wire n_7;
wire n_8;
wire n_9;
wire n_10;
wire n_11;
wire n_12;
wire n_14;
wire n_17;
wire n_19;
wire n_20;
wire n_21;
wire n_22;
wire n_23;
wire n_25;
wire n_26;
wire n_29;
wire n_30;
wire n_32;
wire n_0;
wire n_34;
wire n_33;
wire n_31;
wire slo__sro_n57;
wire slo__sro_n58;
wire slo__sro_n59;
wire slo__sro_n60;
wire slo__sro_n70;
wire slo__sro_n71;
wire slo__sro_n72;
wire slo__sro_n73;
wire slo__sro_n83;
wire slo__sro_n84;
wire slo__sro_n86;
wire slo__sro_n98;
wire slo__sro_n99;
wire slo__sro_n100;
wire slo__sro_n101;
wire slo__sro_n102;
wire slo__sro_n130;
wire slo__sro_n131;
wire slo__sro_n132;
wire slo__sro_n133;
wire slo__sro_n134;
wire slo__sro_n148;
wire slo__sro_n149;
wire slo__sro_n150;
wire slo__sro_n164;
wire slo__sro_n165;
wire slo__sro_n166;
wire slo__sro_n167;
wire slo__sro_n285;
wire slo__sro_n286;
wire slo__sro_n287;
wire slo__sro_n288;
wire slo__sro_n289;
wire slo__sro_n302;
wire slo__sro_n303;
wire slo__sro_n304;
wire slo__sro_n305;
wire slo__sro_n306;
wire slo__sro_n321;
wire slo__sro_n214;
wire slo__sro_n215;
wire slo__sro_n216;
wire slo__sro_n217;
wire slo__sro_n218;
wire slo__sro_n323;
wire slo__sro_n324;
wire slo__sro_n786;
wire slo__sro_n787;
wire slo__sro_n788;
wire slo__sro_n789;
wire slo__n973;
wire slo__sro_n1068;
wire slo__sro_n1069;
wire slo__sro_n1070;
wire slo__sro_n1071;
wire CLOCK_slo__sro_n1150;
wire CLOCK_slo__sro_n1151;
wire CLOCK_slo__sro_n1152;
wire CLOCK_slo__mro_n1241;
wire CLOCK_slo__sro_n1253;
wire CLOCK_slo__sro_n1254;
wire CLOCK_slo__sro_n1255;
wire CLOCK_slo__sro_n1497;
wire CLOCK_slo__sro_n1498;
wire CLOCK_slo__sro_n1499;
wire CLOCK_slo__sro_n1500;
wire CLOCK_slo__mro_n1646;
wire CLOCK_slo__mro_n1645;


INV_X1 i_36 (.ZN (n_34), .A (Multiplier[30]));
INV_X1 i_35 (.ZN (n_33), .A (p_0[30]));
INV_X1 i_34 (.ZN (n_32), .A (n_30));
OAI33_X1 i_33 (.ZN (n_31), .A1 (n_32), .A2 (p_0[30]), .A3 (n_34), .B1 (n_30), .B2 (n_33), .B3 (Multiplier[30]));
XOR2_X1 i_32 (.Z (p_1[31]), .A (Multiplier[31]), .B (n_31));
OAI22_X1 i_31 (.ZN (n_0), .A1 (n_34), .A2 (p_0[30]), .B1 (Multiplier[30]), .B2 (n_33));
XNOR2_X1 i_0 (.ZN (p_1[30]), .A (n_32), .B (n_0));
FA_X1 i_30 (.CO (n_30), .S (p_1[29]), .A (Multiplier[29]), .B (p_0[29]), .CI (n_29));
INV_X1 slo__sro_c98 (.ZN (slo__sro_n167), .A (n_19));
INV_X1 slo__sro_c82 (.ZN (slo__sro_n150), .A (p_0[28]));
INV_X1 slo__sro_c41 (.ZN (slo__sro_n102), .A (n_23));
INV_X1 slo__sro_c15 (.ZN (slo__sro_n73), .A (n_20));
FA_X1 i_25 (.CO (n_25), .S (p_1[24]), .A (Multiplier[24]), .B (p_0[24]), .CI (slo__sro_n99));
INV_X1 slo__sro_c68 (.ZN (slo__sro_n134), .A (p_0[27]));
OAI21_X1 slo__c693 (.ZN (slo__n973), .A (slo__sro_n59), .B1 (slo__sro_n60), .B2 (slo__sro_n58));
FA_X1 i_22 (.CO (n_22), .S (p_1[21]), .A (Multiplier[21]), .B (p_0[21]), .CI (n_21));
NAND2_X1 slo__sro_c29 (.ZN (slo__sro_n86), .A1 (n_26), .A2 (Multiplier[26]));
INV_X1 slo__sro_c212 (.ZN (slo__sro_n289), .A (n_17));
FA_X1 i_19 (.CO (n_19), .S (p_1[18]), .A (Multiplier[18]), .B (p_0[18]), .CI (slo__sro_n286));
INV_X1 slo__sro_c226 (.ZN (slo__sro_n306), .A (n_14));
FA_X1 i_17 (.CO (n_17), .S (p_1[16]), .A (Multiplier[16]), .B (p_0[16]), .CI (slo__sro_n1069));
NAND2_X1 CLOCK_slo__sro_c786 (.ZN (CLOCK_slo__sro_n1152), .A1 (n_4), .A2 (Multiplier[4]));
INV_X1 slo__sro_c242 (.ZN (slo__sro_n324), .A (p_0[13]));
INV_X2 slo__sro_c523 (.ZN (slo__sro_n789), .A (n_22));
NOR2_X1 slo__sro_c244 (.ZN (slo__sro_n322), .A1 (slo__sro_n215), .A2 (Multiplier[13]));
FA_X1 i_12 (.CO (n_12), .S (p_1[11]), .A (Multiplier[11]), .B (p_0[11]), .CI (n_11));
INV_X1 CLOCK_slo__sro_c1112 (.ZN (CLOCK_slo__sro_n1500), .A (p_0[1]));
FA_X1 i_10 (.CO (n_10), .S (p_1[9]), .A (Multiplier[9]), .B (p_0[9]), .CI (n_9));
FA_X1 i_9 (.CO (n_9), .S (p_1[8]), .A (Multiplier[8]), .B (p_0[8]), .CI (n_8));
FA_X1 i_8 (.CO (n_8), .S (p_1[7]), .A (Multiplier[7]), .B (p_0[7]), .CI (n_7));
FA_X1 i_7 (.CO (n_7), .S (p_1[6]), .A (Multiplier[6]), .B (p_0[6]), .CI (n_6));
FA_X1 i_6 (.CO (n_6), .S (p_1[5]), .A (Multiplier[5]), .B (p_0[5]), .CI (n_5));
XNOR2_X2 CLOCK_slo__mro_c884 (.ZN (CLOCK_slo__mro_n1241), .A (slo__sro_n131), .B (Multiplier[28]));
FA_X1 i_4 (.CO (n_4), .S (p_1[3]), .A (Multiplier[3]), .B (p_0[3]), .CI (n_3));
FA_X1 i_3 (.CO (n_3), .S (p_1[2]), .A (Multiplier[2]), .B (p_0[2]), .CI (n_2));
INV_X1 CLOCK_slo__mro_c1244 (.ZN (CLOCK_slo__mro_n1646), .A (p_0[26]));
HA_X1 i_1 (.CO (n_1), .S (p_1[0]), .A (Multiplier[0]), .B (p_0[0]));
INV_X1 slo__sro_c1 (.ZN (slo__sro_n60), .A (n_25));
NAND2_X1 slo__sro_c2 (.ZN (slo__sro_n59), .A1 (p_0[25]), .A2 (Multiplier[25]));
NOR2_X1 slo__sro_c3 (.ZN (slo__sro_n58), .A1 (p_0[25]), .A2 (Multiplier[25]));
OAI21_X1 slo__sro_c4 (.ZN (n_26), .A (slo__sro_n59), .B1 (slo__sro_n58), .B2 (slo__sro_n60));
XNOR2_X2 slo__sro_c5 (.ZN (slo__sro_n57), .A (p_0[25]), .B (Multiplier[25]));
XNOR2_X2 slo__sro_c6 (.ZN (p_1[25]), .A (slo__sro_n57), .B (n_25));
NAND2_X1 slo__sro_c16 (.ZN (slo__sro_n72), .A1 (p_0[20]), .A2 (Multiplier[20]));
NOR2_X1 slo__sro_c17 (.ZN (slo__sro_n71), .A1 (p_0[20]), .A2 (Multiplier[20]));
OAI21_X2 slo__sro_c18 (.ZN (n_21), .A (slo__sro_n72), .B1 (slo__sro_n73), .B2 (slo__sro_n71));
XNOR2_X1 slo__sro_c19 (.ZN (slo__sro_n70), .A (p_0[20]), .B (Multiplier[20]));
XNOR2_X1 slo__sro_c20 (.ZN (p_1[20]), .A (slo__sro_n70), .B (n_20));
XNOR2_X1 slo__sro_c32 (.ZN (slo__sro_n83), .A (slo__n973), .B (Multiplier[26]));
XNOR2_X1 slo__sro_c33 (.ZN (p_1[26]), .A (slo__sro_n83), .B (p_0[26]));
NAND2_X1 slo__sro_c42 (.ZN (slo__sro_n101), .A1 (p_0[23]), .A2 (Multiplier[23]));
NOR2_X1 slo__sro_c43 (.ZN (slo__sro_n100), .A1 (p_0[23]), .A2 (Multiplier[23]));
OAI21_X1 slo__sro_c44 (.ZN (slo__sro_n99), .A (slo__sro_n101), .B1 (slo__sro_n102), .B2 (slo__sro_n100));
XNOR2_X1 slo__sro_c45 (.ZN (slo__sro_n98), .A (p_0[23]), .B (Multiplier[23]));
XNOR2_X1 slo__sro_c46 (.ZN (p_1[23]), .A (slo__sro_n98), .B (n_23));
NAND2_X1 slo__sro_c69 (.ZN (slo__sro_n133), .A1 (slo__sro_n84), .A2 (Multiplier[27]));
NOR2_X2 slo__sro_c70 (.ZN (slo__sro_n132), .A1 (slo__sro_n84), .A2 (Multiplier[27]));
OAI21_X2 slo__sro_c71 (.ZN (slo__sro_n131), .A (slo__sro_n133), .B1 (slo__sro_n132), .B2 (slo__sro_n134));
XNOR2_X1 slo__sro_c72 (.ZN (slo__sro_n130), .A (slo__sro_n84), .B (Multiplier[27]));
XNOR2_X1 slo__sro_c73 (.ZN (p_1[27]), .A (slo__sro_n130), .B (p_0[27]));
NAND2_X1 slo__sro_c83 (.ZN (slo__sro_n149), .A1 (slo__sro_n131), .A2 (Multiplier[28]));
NOR2_X1 slo__sro_c84 (.ZN (slo__sro_n148), .A1 (slo__sro_n131), .A2 (Multiplier[28]));
OAI21_X2 slo__sro_c85 (.ZN (n_29), .A (slo__sro_n149), .B1 (slo__sro_n150), .B2 (slo__sro_n148));
INV_X1 CLOCK_slo__sro_c892 (.ZN (CLOCK_slo__sro_n1255), .A (n_10));
NAND2_X1 CLOCK_slo__sro_c893 (.ZN (CLOCK_slo__sro_n1254), .A1 (p_0[10]), .A2 (Multiplier[10]));
NAND2_X1 slo__sro_c99 (.ZN (slo__sro_n166), .A1 (p_0[19]), .A2 (Multiplier[19]));
NOR2_X1 slo__sro_c100 (.ZN (slo__sro_n165), .A1 (p_0[19]), .A2 (Multiplier[19]));
OAI21_X2 slo__sro_c101 (.ZN (n_20), .A (slo__sro_n166), .B1 (slo__sro_n167), .B2 (slo__sro_n165));
XNOR2_X1 slo__sro_c102 (.ZN (slo__sro_n164), .A (p_0[19]), .B (Multiplier[19]));
XNOR2_X1 slo__sro_c103 (.ZN (p_1[19]), .A (slo__sro_n164), .B (n_19));
NAND2_X1 slo__sro_c213 (.ZN (slo__sro_n288), .A1 (p_0[17]), .A2 (Multiplier[17]));
NOR2_X1 slo__sro_c214 (.ZN (slo__sro_n287), .A1 (p_0[17]), .A2 (Multiplier[17]));
OAI21_X1 slo__sro_c215 (.ZN (slo__sro_n286), .A (slo__sro_n288), .B1 (slo__sro_n289), .B2 (slo__sro_n287));
XNOR2_X1 slo__sro_c216 (.ZN (slo__sro_n285), .A (p_0[17]), .B (Multiplier[17]));
XNOR2_X1 slo__sro_c217 (.ZN (p_1[17]), .A (slo__sro_n285), .B (n_17));
NAND2_X1 slo__sro_c227 (.ZN (slo__sro_n305), .A1 (p_0[14]), .A2 (Multiplier[14]));
NOR2_X2 slo__sro_c228 (.ZN (slo__sro_n304), .A1 (p_0[14]), .A2 (Multiplier[14]));
OAI21_X2 slo__sro_c229 (.ZN (slo__sro_n303), .A (slo__sro_n305), .B1 (slo__sro_n304), .B2 (slo__sro_n306));
XNOR2_X1 slo__sro_c230 (.ZN (slo__sro_n302), .A (p_0[14]), .B (Multiplier[14]));
XNOR2_X1 slo__sro_c231 (.ZN (p_1[14]), .A (slo__sro_n302), .B (n_14));
NAND2_X1 slo__sro_c243 (.ZN (slo__sro_n323), .A1 (slo__sro_n215), .A2 (Multiplier[13]));
INV_X2 slo__sro_c146 (.ZN (slo__sro_n218), .A (n_12));
NAND2_X1 slo__sro_c147 (.ZN (slo__sro_n217), .A1 (p_0[12]), .A2 (Multiplier[12]));
NOR2_X1 slo__sro_c148 (.ZN (slo__sro_n216), .A1 (p_0[12]), .A2 (Multiplier[12]));
OAI21_X2 slo__sro_c149 (.ZN (slo__sro_n215), .A (slo__sro_n217), .B1 (slo__sro_n218), .B2 (slo__sro_n216));
XNOR2_X2 slo__sro_c150 (.ZN (slo__sro_n214), .A (p_0[12]), .B (Multiplier[12]));
XNOR2_X1 slo__sro_c151 (.ZN (p_1[12]), .A (n_12), .B (slo__sro_n214));
OAI21_X2 slo__sro_c245 (.ZN (n_14), .A (slo__sro_n323), .B1 (slo__sro_n322), .B2 (slo__sro_n324));
XNOR2_X2 slo__sro_c246 (.ZN (slo__sro_n321), .A (slo__sro_n215), .B (Multiplier[13]));
XNOR2_X2 slo__sro_c247 (.ZN (p_1[13]), .A (slo__sro_n321), .B (p_0[13]));
NAND2_X1 slo__sro_c524 (.ZN (slo__sro_n788), .A1 (p_0[22]), .A2 (Multiplier[22]));
NOR2_X2 slo__sro_c525 (.ZN (slo__sro_n787), .A1 (p_0[22]), .A2 (Multiplier[22]));
OAI21_X2 slo__sro_c526 (.ZN (n_23), .A (slo__sro_n788), .B1 (slo__sro_n789), .B2 (slo__sro_n787));
XNOR2_X1 slo__sro_c527 (.ZN (slo__sro_n786), .A (p_0[22]), .B (Multiplier[22]));
XNOR2_X1 slo__sro_c528 (.ZN (p_1[22]), .A (slo__sro_n786), .B (n_22));
NAND2_X1 slo__sro_c746 (.ZN (slo__sro_n1071), .A1 (p_0[15]), .A2 (Multiplier[15]));
OAI21_X1 slo__sro_c747 (.ZN (slo__sro_n1070), .A (slo__sro_n303), .B1 (p_0[15]), .B2 (Multiplier[15]));
NAND2_X1 slo__sro_c748 (.ZN (slo__sro_n1069), .A1 (slo__sro_n1070), .A2 (slo__sro_n1071));
XNOR2_X2 slo__sro_c749 (.ZN (slo__sro_n1068), .A (slo__sro_n303), .B (Multiplier[15]));
XNOR2_X2 slo__sro_c750 (.ZN (p_1[15]), .A (slo__sro_n1068), .B (p_0[15]));
OAI21_X1 CLOCK_slo__sro_c787 (.ZN (CLOCK_slo__sro_n1151), .A (p_0[4]), .B1 (n_4), .B2 (Multiplier[4]));
NAND2_X1 CLOCK_slo__sro_c788 (.ZN (n_5), .A1 (CLOCK_slo__sro_n1151), .A2 (CLOCK_slo__sro_n1152));
XNOR2_X2 CLOCK_slo__sro_c789 (.ZN (CLOCK_slo__sro_n1150), .A (n_4), .B (Multiplier[4]));
XNOR2_X2 CLOCK_slo__sro_c790 (.ZN (p_1[4]), .A (CLOCK_slo__sro_n1150), .B (p_0[4]));
XNOR2_X2 CLOCK_slo__mro_c885 (.ZN (p_1[28]), .A (CLOCK_slo__mro_n1241), .B (p_0[28]));
NOR2_X1 CLOCK_slo__sro_c894 (.ZN (CLOCK_slo__sro_n1253), .A1 (p_0[10]), .A2 (Multiplier[10]));
OAI21_X2 CLOCK_slo__sro_c895 (.ZN (n_11), .A (CLOCK_slo__sro_n1254), .B1 (CLOCK_slo__sro_n1255), .B2 (CLOCK_slo__sro_n1253));
XNOR2_X1 CLOCK_slo__sro_c896 (.ZN (CLOCK_slo__sro_n1252), .A (p_0[10]), .B (Multiplier[10]));
XNOR2_X1 CLOCK_slo__sro_c897 (.ZN (p_1[10]), .A (CLOCK_slo__sro_n1252), .B (n_10));
NAND2_X1 CLOCK_slo__sro_c1113 (.ZN (CLOCK_slo__sro_n1499), .A1 (n_1), .A2 (Multiplier[1]));
NOR2_X1 CLOCK_slo__sro_c1114 (.ZN (CLOCK_slo__sro_n1498), .A1 (n_1), .A2 (Multiplier[1]));
OAI21_X1 CLOCK_slo__sro_c1115 (.ZN (n_2), .A (CLOCK_slo__sro_n1499), .B1 (CLOCK_slo__sro_n1500), .B2 (CLOCK_slo__sro_n1498));
XNOR2_X1 CLOCK_slo__sro_c1116 (.ZN (CLOCK_slo__sro_n1497), .A (n_1), .B (Multiplier[1]));
XNOR2_X1 CLOCK_slo__sro_c1117 (.ZN (p_1[1]), .A (CLOCK_slo__sro_n1497), .B (p_0[1]));
NOR2_X2 CLOCK_slo__mro_c1245 (.ZN (CLOCK_slo__mro_n1645), .A1 (n_26), .A2 (Multiplier[26]));
OAI21_X2 CLOCK_slo__mro_c1246 (.ZN (slo__sro_n84), .A (slo__sro_n86), .B1 (CLOCK_slo__mro_n1645), .B2 (CLOCK_slo__mro_n1646));

endmodule //datapath__0_136

module datapath__0_132 (p_1_3_PP_0, p_0, p_1, p_2);

output [31:0] p_2;
input [31:0] p_0;
input [31:0] p_1;
input p_1_3_PP_0;
wire CLOCK_sgo__n1049;
wire CLOCK_slo__sro_n1175;
wire slo__sro_n631;
wire CLOCK_slo__sro_n1395;
wire slo__sro_n630;
wire CLOCK_slo__sro_n1099;
wire n_1;
wire n_2;
wire n_5;
wire n_6;
wire n_8;
wire n_9;
wire n_10;
wire n_11;
wire n_13;
wire n_14;
wire n_15;
wire n_16;
wire n_18;
wire n_19;
wire n_20;
wire n_21;
wire n_23;
wire n_24;
wire n_25;
wire n_26;
wire n_28;
wire n_29;
wire n_30;
wire n_32;
wire n_0;
wire n_34;
wire n_33;
wire n_31;
wire slo__sro_n78;
wire slo__sro_n79;
wire slo__sro_n80;
wire slo__sro_n81;
wire slo__sro_n82;
wire slo__sro_n96;
wire slo__sro_n97;
wire slo__sro_n98;
wire slo__sro_n154;
wire slo__sro_n155;
wire slo__sro_n156;
wire slo__sro_n168;
wire slo__sro_n169;
wire slo__sro_n170;
wire slo__sro_n171;
wire slo__sro_n266;
wire slo__sro_n267;
wire slo__sro_n268;
wire slo__sro_n269;
wire slo__sro_n284;
wire slo__sro_n285;
wire slo__sro_n286;
wire slo__sro_n287;
wire slo__sro_n333;
wire slo__sro_n334;
wire slo__sro_n335;
wire slo__sro_n336;
wire slo__sro_n512;
wire slo__n356;
wire slo__sro_n629;
wire slo__sro_n513;
wire slo__sro_n514;
wire slo__sro_n515;
wire slo__sro_n516;
wire slo__sro_n632;
wire slo__sro_n633;
wire slo__sro_n657;
wire slo__sro_n658;
wire slo__sro_n659;
wire slo__sro_n660;
wire slo__sro_n661;
wire CLOCK_sgo__n1050;
wire CLOCK_slo__mro_n1068;
wire CLOCK_slo__sro_n1100;
wire CLOCK_slo__sro_n1101;
wire CLOCK_slo__sro_n1102;
wire CLOCK_slo__sro_n1114;
wire CLOCK_slo__sro_n1115;
wire CLOCK_slo__sro_n1116;
wire CLOCK_slo__sro_n1117;
wire CLOCK_slo__mro_n1153;
wire CLOCK_slo__sro_n1176;
wire CLOCK_slo__sro_n1177;
wire CLOCK_slo__sro_n1178;
wire CLOCK_slo__mro_n1545;
wire CLOCK_slo__sro_n1396;
wire CLOCK_slo__sro_n1397;
wire CLOCK_slo__sro_n1398;
wire CLOCK_slo__sro_n1221;
wire CLOCK_slo__sro_n1222;
wire CLOCK_slo__sro_n1223;
wire CLOCK_slo__sro_n1224;
wire CLOCK_slo__sro_n1225;
wire CLOCK_slo__sro_n1502;
wire CLOCK_slo__sro_n1503;
wire CLOCK_slo__sro_n1504;
wire CLOCK_slo__sro_n1505;


INV_X1 i_36 (.ZN (n_34), .A (p_0[30]));
INV_X1 i_35 (.ZN (n_33), .A (p_1[30]));
INV_X1 i_34 (.ZN (n_32), .A (n_30));
OAI33_X1 i_33 (.ZN (n_31), .A1 (n_34), .A2 (p_1[30]), .A3 (n_32), .B1 (n_30), .B2 (n_33), .B3 (p_0[30]));
XOR2_X1 i_32 (.Z (p_2[31]), .A (p_0[31]), .B (n_31));
OAI22_X1 i_31 (.ZN (n_0), .A1 (n_34), .A2 (p_1[30]), .B1 (p_0[30]), .B2 (n_33));
XNOR2_X1 i_0 (.ZN (p_2[30]), .A (n_32), .B (n_0));
XNOR2_X1 CLOCK_slo__mro_c717 (.ZN (CLOCK_slo__mro_n1153), .A (p_1[16]), .B (p_0[16]));
FA_X1 i_29 (.CO (n_29), .S (p_2[28]), .A (p_0[28]), .B (p_1[28]), .CI (n_28));
FA_X1 i_28 (.CO (n_28), .S (p_2[27]), .A (p_0[27]), .B (p_1[27]), .CI (slo__sro_n658));
XNOR2_X1 CLOCK_slo__mro_c1051 (.ZN (CLOCK_slo__mro_n1545), .A (p_1[23]), .B (p_0[23]));
FA_X1 i_26 (.CO (n_26), .S (p_2[25]), .A (p_0[25]), .B (p_1[25]), .CI (n_25));
FA_X1 i_25 (.CO (n_25), .S (p_2[24]), .A (p_0[24]), .B (p_1[24]), .CI (n_24));
INV_X1 slo__sro_c97 (.ZN (slo__sro_n171), .A (slo__sro_n513));
INV_X1 slo__sro_c189 (.ZN (slo__sro_n269), .A (n_16));
OAI21_X1 slo__sro_c408 (.ZN (slo__sro_n630), .A (slo__sro_n632), .B1 (slo__sro_n631), .B2 (slo__sro_n633));
FA_X1 i_21 (.CO (n_21), .S (p_2[20]), .A (p_0[20]), .B (p_1[20]), .CI (n_20));
INV_X1 CLOCK_slo__sro_c913 (.ZN (CLOCK_slo__sro_n1398), .A (p_1[1]));
FA_X1 i_19 (.CO (n_19), .S (p_2[18]), .A (p_0[18]), .B (p_1[18]), .CI (n_18));
FA_X1 i_18 (.CO (n_18), .S (p_2[17]), .A (p_0[17]), .B (p_1[17]), .CI (slo__sro_n266));
INV_X1 slo__sro_c205 (.ZN (slo__sro_n287), .A (n_15));
NAND2_X1 slo__sro_c356 (.ZN (slo__sro_n515), .A1 (p_1[21]), .A2 (p_0[21]));
FA_X1 i_15 (.CO (n_15), .S (p_2[14]), .A (p_0[14]), .B (p_1[14]), .CI (n_14));
FA_X1 i_13 (.CO (n_13), .S (p_2[12]), .A (p_0[12]), .B (p_1[12]), .CI (CLOCK_slo__sro_n1222));
NAND2_X1 CLOCK_slo__sro_c1008 (.ZN (CLOCK_slo__sro_n1504), .A1 (p_1[13]), .A2 (p_0[13]));
FA_X1 i_11 (.CO (n_11), .S (p_2[10]), .A (p_0[10]), .B (p_1[10]), .CI (n_10));
FA_X1 i_10 (.CO (n_10), .S (p_2[9]), .A (p_0[9]), .B (p_1[9]), .CI (n_9));
FA_X1 i_9 (.CO (n_9), .S (p_2[8]), .A (p_0[8]), .B (p_1[8]), .CI (n_8));
FA_X1 i_8 (.CO (n_8), .S (p_2[7]), .A (p_0[7]), .B (p_1[7]), .CI (slo__sro_n630));
INV_X1 slo__sro_c428 (.ZN (slo__sro_n661), .A (n_26));
INV_X2 CLOCK_slo__sro_c681 (.ZN (CLOCK_slo__sro_n1117), .A (n_29));
INV_X1 slo__sro_c81 (.ZN (slo__sro_n156), .A (n_23));
NOR2_X1 slo__sro_c407 (.ZN (slo__sro_n631), .A1 (n_6), .A2 (p_0[6]));
INV_X1 slo__sro_c28 (.ZN (slo__sro_n98), .A (slo__sro_n334));
HA_X1 i_1 (.CO (n_1), .S (p_2[0]), .A (p_0[0]), .B (p_1[0]));
INV_X1 slo__sro_c14 (.ZN (slo__sro_n82), .A (n_2));
NAND2_X1 slo__sro_c15 (.ZN (slo__sro_n81), .A1 (p_1[2]), .A2 (p_0[2]));
NOR2_X2 slo__sro_c16 (.ZN (slo__sro_n80), .A1 (p_1[2]), .A2 (p_0[2]));
OAI21_X1 slo__sro_c17 (.ZN (slo__sro_n79), .A (slo__sro_n81), .B1 (slo__sro_n82), .B2 (slo__sro_n80));
XNOR2_X2 slo__sro_c18 (.ZN (slo__sro_n78), .A (p_1[2]), .B (p_0[2]));
XNOR2_X2 slo__sro_c19 (.ZN (p_2[2]), .A (slo__sro_n78), .B (n_2));
NAND2_X1 slo__sro_c29 (.ZN (slo__sro_n97), .A1 (p_1[4]), .A2 (p_0[4]));
NOR2_X1 slo__sro_c30 (.ZN (slo__sro_n96), .A1 (p_1[4]), .A2 (p_0[4]));
OAI21_X1 slo__sro_c31 (.ZN (n_5), .A (slo__sro_n97), .B1 (slo__sro_n96), .B2 (slo__sro_n98));
INV_X1 CLOCK_slo__sro_c665 (.ZN (CLOCK_slo__sro_n1102), .A (n_5));
NAND2_X1 CLOCK_slo__sro_c666 (.ZN (CLOCK_slo__sro_n1101), .A1 (p_1[5]), .A2 (p_0[5]));
NAND2_X1 slo__sro_c82 (.ZN (slo__sro_n155), .A1 (p_1[23]), .A2 (p_0[23]));
NOR2_X1 slo__sro_c83 (.ZN (slo__sro_n154), .A1 (p_1[23]), .A2 (p_0[23]));
OAI21_X1 slo__sro_c84 (.ZN (n_24), .A (slo__sro_n155), .B1 (slo__sro_n156), .B2 (slo__sro_n154));
NAND2_X1 slo__sro_c98 (.ZN (slo__sro_n170), .A1 (p_1[22]), .A2 (p_0[22]));
NOR2_X1 slo__sro_c99 (.ZN (slo__sro_n169), .A1 (p_1[22]), .A2 (p_0[22]));
OAI21_X2 slo__sro_c100 (.ZN (n_23), .A (slo__sro_n170), .B1 (slo__sro_n171), .B2 (slo__sro_n169));
XNOR2_X1 slo__sro_c101 (.ZN (slo__sro_n168), .A (p_1[22]), .B (p_0[22]));
XNOR2_X1 slo__sro_c102 (.ZN (p_2[22]), .A (slo__sro_n168), .B (slo__sro_n513));
NAND2_X1 slo__sro_c190 (.ZN (slo__sro_n268), .A1 (p_1[16]), .A2 (p_0[16]));
NOR2_X1 slo__sro_c191 (.ZN (slo__sro_n267), .A1 (p_1[16]), .A2 (p_0[16]));
OAI21_X2 slo__sro_c192 (.ZN (slo__sro_n266), .A (slo__sro_n268), .B1 (slo__sro_n269), .B2 (slo__sro_n267));
INV_X1 CLOCK_slo__sro_c739 (.ZN (CLOCK_slo__sro_n1178), .A (n_19));
NAND2_X1 CLOCK_slo__sro_c740 (.ZN (CLOCK_slo__sro_n1177), .A1 (p_1[19]), .A2 (p_0[19]));
NAND2_X1 slo__sro_c206 (.ZN (slo__sro_n286), .A1 (p_1[15]), .A2 (p_0[15]));
NOR2_X1 slo__sro_c207 (.ZN (slo__sro_n285), .A1 (p_1[15]), .A2 (p_0[15]));
OAI21_X2 slo__sro_c208 (.ZN (n_16), .A (slo__sro_n286), .B1 (slo__sro_n287), .B2 (slo__sro_n285));
XNOR2_X1 slo__sro_c209 (.ZN (slo__sro_n284), .A (p_1[15]), .B (p_0[15]));
XNOR2_X1 slo__sro_c210 (.ZN (p_2[15]), .A (slo__sro_n284), .B (n_15));
XNOR2_X2 CLOCK_slo__mro_c639 (.ZN (CLOCK_slo__mro_n1068), .A (slo__sro_n334), .B (p_0[4]));
NAND2_X1 slo__sro_c232 (.ZN (slo__sro_n336), .A1 (slo__sro_n79), .A2 (p_0[3]));
NOR2_X1 slo__sro_c233 (.ZN (slo__sro_n335), .A1 (slo__sro_n79), .A2 (p_0[3]));
OAI21_X4 slo__sro_c234 (.ZN (slo__sro_n334), .A (slo__sro_n336), .B1 (CLOCK_sgo__n1049), .B2 (slo__sro_n335));
XNOR2_X1 slo__sro_c235 (.ZN (slo__sro_n333), .A (slo__n356), .B (p_0[3]));
XNOR2_X1 slo__sro_c236 (.ZN (p_2[3]), .A (p_1[3]), .B (slo__sro_n333));
INV_X1 slo__sro_c355 (.ZN (slo__sro_n516), .A (n_21));
OAI21_X1 slo__c251 (.ZN (slo__n356), .A (slo__sro_n81), .B1 (slo__sro_n82), .B2 (slo__sro_n80));
NAND2_X1 slo__sro_c406 (.ZN (slo__sro_n632), .A1 (n_6), .A2 (p_0[6]));
INV_X1 slo__sro_c405 (.ZN (slo__sro_n633), .A (p_1[6]));
NOR2_X1 slo__sro_c357 (.ZN (slo__sro_n514), .A1 (p_1[21]), .A2 (p_0[21]));
OAI21_X2 slo__sro_c358 (.ZN (slo__sro_n513), .A (slo__sro_n515), .B1 (slo__sro_n516), .B2 (slo__sro_n514));
XNOR2_X1 slo__sro_c359 (.ZN (slo__sro_n512), .A (p_1[21]), .B (p_0[21]));
XNOR2_X1 slo__sro_c360 (.ZN (p_2[21]), .A (n_21), .B (slo__sro_n512));
XNOR2_X1 slo__sro_c409 (.ZN (slo__sro_n629), .A (n_6), .B (p_0[6]));
XNOR2_X1 slo__sro_c410 (.ZN (p_2[6]), .A (slo__sro_n629), .B (p_1[6]));
NAND2_X1 slo__sro_c429 (.ZN (slo__sro_n660), .A1 (p_1[26]), .A2 (p_0[26]));
NOR2_X1 slo__sro_c430 (.ZN (slo__sro_n659), .A1 (p_1[26]), .A2 (p_0[26]));
OAI21_X2 slo__sro_c431 (.ZN (slo__sro_n658), .A (slo__sro_n660), .B1 (slo__sro_n661), .B2 (slo__sro_n659));
XNOR2_X2 slo__sro_c432 (.ZN (slo__sro_n657), .A (p_1[26]), .B (p_0[26]));
XNOR2_X2 slo__sro_c433 (.ZN (p_2[26]), .A (slo__sro_n657), .B (n_26));
INV_X2 CLOCK_sgo__L3_c5_c631 (.ZN (CLOCK_sgo__n1049), .A (CLOCK_sgo__n1050));
BUF_X1 CLOCK_sgo__L2_c4_c632 (.Z (CLOCK_sgo__n1050), .A (p_1_3_PP_0));
XNOR2_X2 CLOCK_slo__mro_c640 (.ZN (p_2[4]), .A (CLOCK_slo__mro_n1068), .B (p_1[4]));
NOR2_X1 CLOCK_slo__sro_c667 (.ZN (CLOCK_slo__sro_n1100), .A1 (p_1[5]), .A2 (p_0[5]));
OAI21_X2 CLOCK_slo__sro_c668 (.ZN (n_6), .A (CLOCK_slo__sro_n1101), .B1 (CLOCK_slo__sro_n1102), .B2 (CLOCK_slo__sro_n1100));
XNOR2_X2 CLOCK_slo__sro_c669 (.ZN (CLOCK_slo__sro_n1099), .A (p_1[5]), .B (p_0[5]));
XNOR2_X2 CLOCK_slo__sro_c670 (.ZN (p_2[5]), .A (CLOCK_slo__sro_n1099), .B (n_5));
NAND2_X1 CLOCK_slo__sro_c682 (.ZN (CLOCK_slo__sro_n1116), .A1 (p_1[29]), .A2 (p_0[29]));
NOR2_X1 CLOCK_slo__sro_c683 (.ZN (CLOCK_slo__sro_n1115), .A1 (p_1[29]), .A2 (p_0[29]));
OAI21_X2 CLOCK_slo__sro_c684 (.ZN (n_30), .A (CLOCK_slo__sro_n1116), .B1 (CLOCK_slo__sro_n1117), .B2 (CLOCK_slo__sro_n1115));
XNOR2_X1 CLOCK_slo__sro_c685 (.ZN (CLOCK_slo__sro_n1114), .A (p_1[29]), .B (p_0[29]));
XNOR2_X1 CLOCK_slo__sro_c686 (.ZN (p_2[29]), .A (n_29), .B (CLOCK_slo__sro_n1114));
XNOR2_X1 CLOCK_slo__mro_c718 (.ZN (p_2[16]), .A (CLOCK_slo__mro_n1153), .B (n_16));
NOR2_X1 CLOCK_slo__sro_c741 (.ZN (CLOCK_slo__sro_n1176), .A1 (p_1[19]), .A2 (p_0[19]));
OAI21_X1 CLOCK_slo__sro_c742 (.ZN (n_20), .A (CLOCK_slo__sro_n1177), .B1 (CLOCK_slo__sro_n1178), .B2 (CLOCK_slo__sro_n1176));
XNOR2_X1 CLOCK_slo__sro_c743 (.ZN (CLOCK_slo__sro_n1175), .A (p_1[19]), .B (p_0[19]));
XNOR2_X1 CLOCK_slo__sro_c744 (.ZN (p_2[19]), .A (CLOCK_slo__sro_n1175), .B (n_19));
XNOR2_X1 CLOCK_slo__mro_c1052 (.ZN (p_2[23]), .A (CLOCK_slo__mro_n1545), .B (n_23));
NAND2_X1 CLOCK_slo__sro_c914 (.ZN (CLOCK_slo__sro_n1397), .A1 (n_1), .A2 (p_0[1]));
NOR2_X1 CLOCK_slo__sro_c915 (.ZN (CLOCK_slo__sro_n1396), .A1 (n_1), .A2 (p_0[1]));
OAI21_X2 CLOCK_slo__sro_c916 (.ZN (n_2), .A (CLOCK_slo__sro_n1397), .B1 (CLOCK_slo__sro_n1396), .B2 (CLOCK_slo__sro_n1398));
XNOR2_X1 CLOCK_slo__sro_c917 (.ZN (CLOCK_slo__sro_n1395), .A (n_1), .B (p_0[1]));
XNOR2_X1 CLOCK_slo__sro_c918 (.ZN (p_2[1]), .A (CLOCK_slo__sro_n1395), .B (p_1[1]));
INV_X1 CLOCK_slo__sro_c1007 (.ZN (CLOCK_slo__sro_n1505), .A (n_13));
INV_X1 CLOCK_slo__sro_c783 (.ZN (CLOCK_slo__sro_n1225), .A (n_11));
NAND2_X1 CLOCK_slo__sro_c784 (.ZN (CLOCK_slo__sro_n1224), .A1 (p_1[11]), .A2 (p_0[11]));
NOR2_X1 CLOCK_slo__sro_c785 (.ZN (CLOCK_slo__sro_n1223), .A1 (p_1[11]), .A2 (p_0[11]));
OAI21_X1 CLOCK_slo__sro_c786 (.ZN (CLOCK_slo__sro_n1222), .A (CLOCK_slo__sro_n1224)
    , .B1 (CLOCK_slo__sro_n1225), .B2 (CLOCK_slo__sro_n1223));
XNOR2_X1 CLOCK_slo__sro_c787 (.ZN (CLOCK_slo__sro_n1221), .A (p_1[11]), .B (p_0[11]));
XNOR2_X1 CLOCK_slo__sro_c788 (.ZN (p_2[11]), .A (n_11), .B (CLOCK_slo__sro_n1221));
NOR2_X1 CLOCK_slo__sro_c1009 (.ZN (CLOCK_slo__sro_n1503), .A1 (p_1[13]), .A2 (p_0[13]));
OAI21_X1 CLOCK_slo__sro_c1010 (.ZN (n_14), .A (CLOCK_slo__sro_n1504), .B1 (CLOCK_slo__sro_n1505), .B2 (CLOCK_slo__sro_n1503));
XNOR2_X1 CLOCK_slo__sro_c1011 (.ZN (CLOCK_slo__sro_n1502), .A (p_1[13]), .B (p_0[13]));
XNOR2_X1 CLOCK_slo__sro_c1012 (.ZN (p_2[13]), .A (n_13), .B (CLOCK_slo__sro_n1502));

endmodule //datapath__0_132

module datapath__0_131 (p_0_1_PP_0, Multiplier, p_0, p_1);

output [31:0] p_1;
input [31:0] Multiplier;
input [31:0] p_0;
input p_0_1_PP_0;
wire CLOCK_slo__xsl_n1785;
wire CLOCK_slo__xsl_n1786;
wire CLOCK_slo__sro_n1328;
wire n_1;
wire CLOCK_slo__sro_n1294;
wire n_3;
wire n_4;
wire n_6;
wire n_7;
wire slo__sro_n868;
wire n_9;
wire n_10;
wire n_11;
wire n_12;
wire n_14;
wire n_15;
wire n_16;
wire n_17;
wire n_18;
wire n_20;
wire slo__xsl_n812;
wire slo__xsl_n824;
wire n_24;
wire slo__sro_n123;
wire n_26;
wire n_27;
wire n_29;
wire n_30;
wire n_32;
wire n_0;
wire n_34;
wire n_33;
wire n_31;
wire slo__sro_n106;
wire slo__sro_n107;
wire slo__sro_n108;
wire slo__sro_n109;
wire slo__sro_n110;
wire slo__sro_n89;
wire slo__sro_n90;
wire slo__sro_n91;
wire slo__sro_n92;
wire slo__sro_n93;
wire slo__sro_n124;
wire slo__sro_n125;
wire slo__sro_n126;
wire slo__sro_n136;
wire slo__sro_n137;
wire slo__sro_n138;
wire slo__sro_n139;
wire slo__sro_n140;
wire slo__sro_n141;
wire slo__sro_n142;
wire slo__sro_n223;
wire slo__sro_n224;
wire slo__sro_n225;
wire slo__sro_n226;
wire slo__sro_n242;
wire slo__sro_n243;
wire slo__sro_n254;
wire slo__sro_n255;
wire slo__sro_n256;
wire slo__sro_n257;
wire slo__sro_n258;
wire slo__xsl_n811;
wire slo__sro_n480;
wire slo__sro_n481;
wire slo__sro_n482;
wire slo__sro_n483;
wire slo__sro_n484;
wire slo__xsl_n825;
wire slo__mro_n853;
wire slo__sro_n869;
wire slo__sro_n870;
wire slo__sro_n871;
wire slo__sro_n872;
wire slo__sro_n933;
wire slo__sro_n934;
wire slo__sro_n935;
wire slo__sro_n936;
wire slo__sro_n937;
wire CLOCK_slo__mro_n1283;
wire CLOCK_slo__sro_n1295;
wire CLOCK_slo__sro_n1296;
wire CLOCK_slo__sro_n1297;
wire CLOCK_slo__sro_n1298;
wire CLOCK_slo__sro_n1315;
wire CLOCK_slo__sro_n1316;
wire CLOCK_slo__sro_n1317;
wire CLOCK_slo__sro_n1318;
wire CLOCK_slo__sro_n1329;
wire CLOCK_slo__sro_n1330;
wire CLOCK_slo__sro_n1331;
wire CLOCK_slo__sro_n1375;
wire CLOCK_slo__sro_n1376;
wire CLOCK_slo__sro_n1377;
wire CLOCK_slo__sro_n1378;
wire CLOCK_slo__sro_n1379;
wire CLOCK_slo__sro_n1392;
wire CLOCK_slo__sro_n1393;
wire CLOCK_slo__sro_n1394;
wire CLOCK_slo__sro_n1395;
wire CLOCK_slo__sro_n1396;
wire CLOCK_slo__sro_n1409;
wire CLOCK_slo__sro_n1410;
wire CLOCK_slo__sro_n1411;
wire CLOCK_slo__sro_n1412;
wire CLOCK_slo__sro_n1715;
wire CLOCK_slo__sro_n1716;
wire CLOCK_slo__sro_n1717;
wire CLOCK_slo__sro_n1718;


INV_X1 i_36 (.ZN (n_34), .A (Multiplier[30]));
INV_X1 i_35 (.ZN (n_33), .A (p_0[30]));
INV_X1 i_34 (.ZN (n_32), .A (n_30));
INV_X2 CLOCK_slo__sro_c983 (.ZN (CLOCK_slo__sro_n1379), .A (n_12));
XOR2_X1 i_32 (.Z (p_1[31]), .A (Multiplier[31]), .B (n_31));
OAI22_X1 i_31 (.ZN (n_0), .A1 (n_34), .A2 (p_0[30]), .B1 (Multiplier[30]), .B2 (n_33));
XNOR2_X1 i_0 (.ZN (p_1[30]), .A (n_32), .B (n_0));
FA_X1 i_30 (.CO (n_30), .S (p_1[29]), .A (Multiplier[29]), .B (p_0[29]), .CI (n_29));
FA_X1 i_29 (.CO (n_29), .S (p_1[28]), .A (Multiplier[28]), .B (p_0[28]), .CI (CLOCK_slo__sro_n1393));
INV_X1 CLOCK_slo__sro_c1011 (.ZN (CLOCK_slo__sro_n1412), .A (n_15));
INV_X1 slo__sro_c71 (.ZN (slo__sro_n142), .A (Multiplier[1]));
INV_X1 CLOCK_slo__xsl_c1337 (.ZN (CLOCK_slo__xsl_n1786), .A (slo__sro_n934));
NAND2_X1 slo__sro_c58 (.ZN (slo__sro_n125), .A1 (p_0[26]), .A2 (Multiplier[26]));
INV_X1 slo__sro_c180 (.ZN (slo__sro_n258), .A (n_20));
INV_X1 slo__sro_c57 (.ZN (slo__sro_n126), .A (n_26));
INV_X1 slo__xsl_c566 (.ZN (slo__xsl_n811), .A (slo__xsl_n812));
INV_X1 slo__xsl_c576 (.ZN (slo__xsl_n825), .A (slo__sro_n481));
INV_X1 CLOCK_slo__sro_c900 (.ZN (CLOCK_slo__sro_n1298), .A (n_4));
FA_X1 i_18 (.CO (n_18), .S (p_1[17]), .A (Multiplier[17]), .B (p_0[17]), .CI (n_17));
FA_X1 i_17 (.CO (n_17), .S (p_1[16]), .A (Multiplier[16]), .B (p_0[16]), .CI (n_16));
INV_X1 CLOCK_slo__sro_c1257 (.ZN (CLOCK_slo__sro_n1718), .A (slo__sro_n934));
FA_X1 i_15 (.CO (n_15), .S (p_1[14]), .A (Multiplier[14]), .B (p_0[14]), .CI (n_14));
FA_X1 i_14 (.CO (n_14), .S (p_1[13]), .A (Multiplier[13]), .B (p_0[13]), .CI (CLOCK_slo__sro_n1376));
NAND2_X1 CLOCK_slo__sro_c997 (.ZN (CLOCK_slo__sro_n1396), .A1 (p_0[27]), .A2 (Multiplier[27]));
FA_X1 i_12 (.CO (n_12), .S (p_1[11]), .A (Multiplier[11]), .B (p_0[11]), .CI (n_11));
FA_X1 i_11 (.CO (n_11), .S (p_1[10]), .A (Multiplier[10]), .B (p_0[10]), .CI (n_10));
FA_X1 i_10 (.CO (n_10), .S (p_1[9]), .A (Multiplier[9]), .B (p_0[9]), .CI (n_9));
INV_X1 CLOCK_slo__sro_c932 (.ZN (CLOCK_slo__sro_n1331), .A (n_30));
NAND2_X1 slo__sro_c168 (.ZN (slo__sro_n243), .A1 (p_0[23]), .A2 (Multiplier[23]));
FA_X1 i_7 (.CO (n_7), .S (p_1[6]), .A (Multiplier[6]), .B (p_0[6]), .CI (n_6));
FA_X1 i_6 (.CO (n_6), .S (p_1[5]), .A (Multiplier[5]), .B (p_0[5]), .CI (CLOCK_slo__sro_n1295));
NAND2_X1 CLOCK_slo__sro_c918 (.ZN (CLOCK_slo__sro_n1318), .A1 (p_0[8]), .A2 (Multiplier[8]));
FA_X1 i_4 (.CO (n_4), .S (p_1[3]), .A (Multiplier[3]), .B (p_0[3]), .CI (n_3));
FA_X1 i_3 (.CO (n_3), .S (p_1[2]), .A (Multiplier[2]), .B (p_0[2]), .CI (slo__sro_n137));
INV_X1 slo__sro_c152 (.ZN (slo__sro_n226), .A (n_7));
HA_X1 i_1 (.CO (n_1), .S (p_1[0]), .A (Multiplier[0]), .B (p_0[0]));
INV_X2 slo__sro_c43 (.ZN (slo__sro_n110), .A (slo__sro_n481));
NAND2_X1 slo__sro_c44 (.ZN (slo__sro_n109), .A1 (p_0[22]), .A2 (Multiplier[22]));
NOR2_X2 slo__sro_c45 (.ZN (slo__sro_n108), .A1 (p_0[22]), .A2 (Multiplier[22]));
OAI21_X1 CLOCK_slo__sro_c1260 (.ZN (n_20), .A (CLOCK_slo__sro_n1717), .B1 (CLOCK_slo__sro_n1716), .B2 (CLOCK_slo__sro_n1718));
XNOR2_X1 slo__sro_c47 (.ZN (slo__sro_n106), .A (p_0[22]), .B (Multiplier[22]));
XNOR2_X2 slo__sro_c48 (.ZN (p_1[22]), .A (slo__sro_n106), .B (slo__xsl_n824));
INV_X1 slo__sro_c29 (.ZN (slo__sro_n93), .A (n_24));
NAND2_X1 slo__sro_c30 (.ZN (slo__sro_n92), .A1 (p_0[24]), .A2 (Multiplier[24]));
NOR2_X1 slo__sro_c31 (.ZN (slo__sro_n91), .A1 (p_0[24]), .A2 (Multiplier[24]));
OAI21_X1 slo__sro_c32 (.ZN (slo__sro_n90), .A (slo__sro_n92), .B1 (slo__sro_n93), .B2 (slo__sro_n91));
XNOR2_X2 slo__sro_c33 (.ZN (slo__sro_n89), .A (p_0[24]), .B (Multiplier[24]));
XNOR2_X2 slo__sro_c34 (.ZN (p_1[24]), .A (slo__sro_n89), .B (n_24));
NOR2_X1 slo__sro_c59 (.ZN (slo__sro_n124), .A1 (p_0[26]), .A2 (Multiplier[26]));
OAI21_X2 slo__sro_c60 (.ZN (n_27), .A (slo__sro_n125), .B1 (slo__sro_n126), .B2 (slo__sro_n124));
XNOR2_X2 slo__sro_c61 (.ZN (slo__sro_n123), .A (p_0[26]), .B (Multiplier[26]));
XNOR2_X2 slo__sro_c62 (.ZN (p_1[26]), .A (slo__sro_n123), .B (n_26));
INV_X1 slo__sro_c72 (.ZN (slo__sro_n141), .A (n_1));
NAND2_X1 slo__sro_c73 (.ZN (slo__sro_n140), .A1 (n_1), .A2 (Multiplier[1]));
NAND2_X2 slo__sro_c74 (.ZN (slo__sro_n139), .A1 (slo__sro_n141), .A2 (slo__sro_n142));
NAND2_X1 slo__sro_c75 (.ZN (slo__sro_n138), .A1 (p_0[1]), .A2 (slo__sro_n139));
NAND2_X2 slo__sro_c76 (.ZN (slo__sro_n137), .A1 (slo__sro_n138), .A2 (slo__sro_n140));
XNOR2_X1 slo__sro_c77 (.ZN (slo__sro_n136), .A (n_1), .B (Multiplier[1]));
XNOR2_X1 slo__sro_c78 (.ZN (p_1[1]), .A (slo__sro_n136), .B (p_0_1_PP_0));
NAND2_X1 slo__sro_c153 (.ZN (slo__sro_n225), .A1 (p_0[7]), .A2 (Multiplier[7]));
NOR2_X1 slo__sro_c154 (.ZN (slo__sro_n224), .A1 (p_0[7]), .A2 (Multiplier[7]));
OAI21_X2 slo__sro_c155 (.ZN (slo__sro_n223), .A (slo__sro_n225), .B1 (slo__sro_n226), .B2 (slo__sro_n224));
XNOR2_X1 CLOCK_slo__mro_c892 (.ZN (CLOCK_slo__mro_n1283), .A (p_0[7]), .B (Multiplier[7]));
NAND2_X1 CLOCK_slo__sro_c901 (.ZN (CLOCK_slo__sro_n1297), .A1 (p_0[4]), .A2 (Multiplier[4]));
AOI22_X1 slo__sro_c169 (.ZN (slo__sro_n242), .A1 (p_0[23]), .A2 (slo__sro_n107), .B1 (slo__sro_n107), .B2 (Multiplier[23]));
NAND2_X1 slo__sro_c170 (.ZN (n_24), .A1 (slo__sro_n243), .A2 (slo__sro_n242));
BUF_X2 slo__sro_c609 (.Z (slo__sro_n872), .A (slo__sro_n90));
NAND2_X1 slo__sro_c610 (.ZN (slo__sro_n871), .A1 (p_0[25]), .A2 (Multiplier[25]));
NAND2_X1 slo__sro_c181 (.ZN (slo__sro_n257), .A1 (p_0[20]), .A2 (Multiplier[20]));
NOR2_X1 slo__sro_c182 (.ZN (slo__sro_n256), .A1 (p_0[20]), .A2 (Multiplier[20]));
OAI21_X2 slo__sro_c183 (.ZN (slo__sro_n255), .A (slo__sro_n257), .B1 (slo__sro_n258), .B2 (slo__sro_n256));
XNOR2_X2 slo__sro_c184 (.ZN (slo__sro_n254), .A (p_0[20]), .B (Multiplier[20]));
XNOR2_X1 slo__sro_c185 (.ZN (p_1[20]), .A (n_20), .B (slo__sro_n254));
INV_X1 slo__xsl_c565 (.ZN (slo__xsl_n812), .A (slo__sro_n255));
INV_X1 slo__sro_c331 (.ZN (slo__sro_n484), .A (slo__sro_n255));
NAND2_X1 slo__sro_c332 (.ZN (slo__sro_n483), .A1 (p_0[21]), .A2 (Multiplier[21]));
NOR2_X2 slo__sro_c333 (.ZN (slo__sro_n482), .A1 (p_0[21]), .A2 (Multiplier[21]));
OAI21_X2 slo__sro_c334 (.ZN (slo__sro_n481), .A (slo__sro_n483), .B1 (slo__sro_n482), .B2 (slo__sro_n484));
XNOR2_X1 slo__sro_c335 (.ZN (slo__sro_n480), .A (p_0[21]), .B (Multiplier[21]));
XNOR2_X1 slo__sro_c336 (.ZN (p_1[21]), .A (slo__sro_n480), .B (slo__xsl_n811));
INV_X1 slo__xsl_c577 (.ZN (slo__xsl_n824), .A (slo__xsl_n825));
XNOR2_X2 slo__mro_c599 (.ZN (slo__mro_n853), .A (slo__sro_n107), .B (Multiplier[23]));
XNOR2_X2 slo__mro_c600 (.ZN (p_1[23]), .A (slo__mro_n853), .B (p_0[23]));
NAND2_X1 slo__sro_c611 (.ZN (slo__sro_n870), .A1 (slo__sro_n872), .A2 (Multiplier[25]));
NAND2_X1 slo__sro_c612 (.ZN (slo__sro_n869), .A1 (slo__sro_n872), .A2 (p_0[25]));
NAND3_X2 slo__sro_c613 (.ZN (n_26), .A1 (slo__sro_n869), .A2 (slo__sro_n870), .A3 (slo__sro_n871));
XNOR2_X2 slo__sro_c614 (.ZN (slo__sro_n868), .A (p_0[25]), .B (Multiplier[25]));
XNOR2_X2 slo__sro_c615 (.ZN (p_1[25]), .A (slo__sro_n868), .B (slo__sro_n872));
INV_X1 CLOCK_slo__xsl_c1338 (.ZN (CLOCK_slo__xsl_n1785), .A (CLOCK_slo__xsl_n1786));
INV_X1 slo__sro_c668 (.ZN (slo__sro_n937), .A (n_18));
NAND2_X1 slo__sro_c669 (.ZN (slo__sro_n936), .A1 (p_0[18]), .A2 (Multiplier[18]));
NOR2_X1 slo__sro_c670 (.ZN (slo__sro_n935), .A1 (p_0[18]), .A2 (Multiplier[18]));
OAI21_X1 slo__sro_c671 (.ZN (slo__sro_n934), .A (slo__sro_n936), .B1 (slo__sro_n937), .B2 (slo__sro_n935));
XNOR2_X1 slo__sro_c672 (.ZN (slo__sro_n933), .A (p_0[18]), .B (Multiplier[18]));
XNOR2_X1 slo__sro_c673 (.ZN (p_1[18]), .A (n_18), .B (slo__sro_n933));
XNOR2_X1 CLOCK_slo__mro_c893 (.ZN (p_1[7]), .A (CLOCK_slo__mro_n1283), .B (n_7));
NOR2_X1 CLOCK_slo__sro_c902 (.ZN (CLOCK_slo__sro_n1296), .A1 (p_0[4]), .A2 (Multiplier[4]));
OAI21_X1 CLOCK_slo__sro_c903 (.ZN (CLOCK_slo__sro_n1295), .A (CLOCK_slo__sro_n1297)
    , .B1 (CLOCK_slo__sro_n1296), .B2 (CLOCK_slo__sro_n1298));
XNOR2_X1 CLOCK_slo__sro_c904 (.ZN (CLOCK_slo__sro_n1294), .A (p_0[4]), .B (Multiplier[4]));
XNOR2_X1 CLOCK_slo__sro_c905 (.ZN (p_1[4]), .A (CLOCK_slo__sro_n1294), .B (n_4));
NAND2_X1 CLOCK_slo__sro_c919 (.ZN (CLOCK_slo__sro_n1317), .A1 (slo__sro_n223), .A2 (Multiplier[8]));
NAND2_X1 CLOCK_slo__sro_c920 (.ZN (CLOCK_slo__sro_n1316), .A1 (slo__sro_n223), .A2 (p_0[8]));
NAND3_X2 CLOCK_slo__sro_c921 (.ZN (n_9), .A1 (CLOCK_slo__sro_n1317), .A2 (CLOCK_slo__sro_n1316), .A3 (CLOCK_slo__sro_n1318));
XNOR2_X2 CLOCK_slo__sro_c922 (.ZN (CLOCK_slo__sro_n1315), .A (p_0[8]), .B (Multiplier[8]));
XNOR2_X2 CLOCK_slo__sro_c923 (.ZN (p_1[8]), .A (CLOCK_slo__sro_n1315), .B (slo__sro_n223));
NOR2_X1 CLOCK_slo__sro_c933 (.ZN (CLOCK_slo__sro_n1330), .A1 (n_33), .A2 (Multiplier[30]));
NAND2_X1 CLOCK_slo__sro_c934 (.ZN (CLOCK_slo__sro_n1329), .A1 (CLOCK_slo__sro_n1330), .A2 (CLOCK_slo__sro_n1331));
OR2_X1 CLOCK_slo__sro_c935 (.ZN (CLOCK_slo__sro_n1328), .A1 (p_0[30]), .A2 (n_34));
OAI21_X1 CLOCK_slo__sro_c936 (.ZN (n_31), .A (CLOCK_slo__sro_n1329), .B1 (n_32), .B2 (CLOCK_slo__sro_n1328));
NAND2_X1 CLOCK_slo__sro_c984 (.ZN (CLOCK_slo__sro_n1378), .A1 (p_0[12]), .A2 (Multiplier[12]));
NOR2_X1 CLOCK_slo__sro_c985 (.ZN (CLOCK_slo__sro_n1377), .A1 (p_0[12]), .A2 (Multiplier[12]));
OAI21_X2 CLOCK_slo__sro_c986 (.ZN (CLOCK_slo__sro_n1376), .A (CLOCK_slo__sro_n1378)
    , .B1 (CLOCK_slo__sro_n1379), .B2 (CLOCK_slo__sro_n1377));
XNOR2_X1 CLOCK_slo__sro_c987 (.ZN (CLOCK_slo__sro_n1375), .A (p_0[12]), .B (Multiplier[12]));
XNOR2_X1 CLOCK_slo__sro_c988 (.ZN (p_1[12]), .A (CLOCK_slo__sro_n1375), .B (n_12));
NAND2_X1 CLOCK_slo__sro_c998 (.ZN (CLOCK_slo__sro_n1395), .A1 (n_27), .A2 (Multiplier[27]));
NAND2_X1 CLOCK_slo__sro_c999 (.ZN (CLOCK_slo__sro_n1394), .A1 (n_27), .A2 (p_0[27]));
NAND3_X1 CLOCK_slo__sro_c1000 (.ZN (CLOCK_slo__sro_n1393), .A1 (CLOCK_slo__sro_n1396)
    , .A2 (CLOCK_slo__sro_n1394), .A3 (CLOCK_slo__sro_n1395));
XNOR2_X1 CLOCK_slo__sro_c1001 (.ZN (CLOCK_slo__sro_n1392), .A (p_0[27]), .B (Multiplier[27]));
XNOR2_X1 CLOCK_slo__sro_c1002 (.ZN (p_1[27]), .A (CLOCK_slo__sro_n1392), .B (n_27));
NAND2_X1 CLOCK_slo__sro_c1012 (.ZN (CLOCK_slo__sro_n1411), .A1 (p_0[15]), .A2 (Multiplier[15]));
NOR2_X1 CLOCK_slo__sro_c1013 (.ZN (CLOCK_slo__sro_n1410), .A1 (p_0[15]), .A2 (Multiplier[15]));
OAI21_X1 CLOCK_slo__sro_c1014 (.ZN (n_16), .A (CLOCK_slo__sro_n1411), .B1 (CLOCK_slo__sro_n1412), .B2 (CLOCK_slo__sro_n1410));
XNOR2_X1 CLOCK_slo__sro_c1015 (.ZN (CLOCK_slo__sro_n1409), .A (p_0[15]), .B (Multiplier[15]));
XNOR2_X1 CLOCK_slo__sro_c1016 (.ZN (p_1[15]), .A (CLOCK_slo__sro_n1409), .B (n_15));
NAND2_X1 CLOCK_slo__sro_c1258 (.ZN (CLOCK_slo__sro_n1717), .A1 (p_0[19]), .A2 (Multiplier[19]));
NOR2_X1 CLOCK_slo__sro_c1259 (.ZN (CLOCK_slo__sro_n1716), .A1 (p_0[19]), .A2 (Multiplier[19]));
OAI21_X2 CLOCK_slo__sro_c1033 (.ZN (slo__sro_n107), .A (slo__sro_n109), .B1 (slo__sro_n110), .B2 (slo__sro_n108));
XNOR2_X1 CLOCK_slo__sro_c1261 (.ZN (CLOCK_slo__sro_n1715), .A (p_0[19]), .B (Multiplier[19]));
XNOR2_X1 CLOCK_slo__sro_c1262 (.ZN (p_1[19]), .A (CLOCK_slo__sro_n1715), .B (CLOCK_slo__xsl_n1785));

endmodule //datapath__0_131

module datapath__0_127 (p_0, p_1, p_2);

output [31:0] p_2;
input [31:0] p_0;
input [31:0] p_1;
wire slo__sro_n775;
wire n_1;
wire slo__sro_n774;
wire n_3;
wire n_4;
wire n_5;
wire n_6;
wire n_7;
wire n_8;
wire n_10;
wire slo__sro_n385;
wire n_13;
wire n_14;
wire n_16;
wire n_18;
wire n_19;
wire n_20;
wire n_21;
wire n_22;
wire n_23;
wire n_27;
wire n_28;
wire n_29;
wire n_30;
wire n_32;
wire n_0;
wire n_34;
wire n_33;
wire n_31;
wire slo__sro_n107;
wire slo__sro_n108;
wire slo__sro_n109;
wire slo__sro_n110;
wire slo__sro_n111;
wire slo__sro_n164;
wire CLOCK_slo__sro_n1109;
wire slo__sro_n166;
wire slo__sro_n167;
wire slo__sro_n268;
wire slo__sro_n269;
wire slo__sro_n270;
wire slo__sro_n271;
wire slo__sro_n272;
wire slo__sro_n285;
wire slo__sro_n286;
wire slo__sro_n287;
wire slo__sro_n288;
wire slo__sro_n289;
wire slo__sro_n302;
wire slo__sro_n303;
wire slo__sro_n304;
wire slo__sro_n305;
wire slo__sro_n306;
wire slo__sro_n383;
wire slo__sro_n384;
wire slo__sro_n251;
wire slo__sro_n252;
wire slo__sro_n253;
wire slo__sro_n254;
wire slo__sro_n255;
wire slo__sro_n386;
wire slo__sro_n601;
wire slo__sro_n423;
wire slo__sro_n424;
wire slo__sro_n425;
wire slo__sro_n426;
wire slo__sro_n602;
wire slo__sro_n603;
wire slo__sro_n604;
wire slo__sro_n605;
wire slo__sro_n776;
wire slo__sro_n777;
wire slo__sro_n778;
wire slo__sro_n723;
wire slo__sro_n724;
wire slo__sro_n725;
wire slo__sro_n726;
wire slo__mro_n761;
wire CLOCK_slo__sro_n997;
wire CLOCK_slo__sro_n998;
wire CLOCK_slo__sro_n1010;
wire CLOCK_slo__sro_n1011;
wire CLOCK_slo__sro_n1012;
wire CLOCK_slo__mro_n1049;
wire CLOCK_slo__sro_n1110;
wire CLOCK_slo__sro_n1111;
wire CLOCK_slo__sro_n1112;
wire CLOCK_slo__sro_n1113;
wire CLOCK_slo__sro_n1145;
wire CLOCK_slo__sro_n1146;
wire CLOCK_slo__sro_n1147;
wire CLOCK_slo__sro_n1148;


INV_X1 i_36 (.ZN (n_34), .A (p_0[30]));
INV_X1 i_35 (.ZN (n_33), .A (p_1[30]));
INV_X1 i_34 (.ZN (n_32), .A (n_30));
INV_X2 CLOCK_slo__sro_c678 (.ZN (CLOCK_slo__sro_n997), .A (p_1[0]));
XOR2_X1 i_32 (.Z (p_2[31]), .A (p_0[31]), .B (n_31));
OAI22_X1 i_31 (.ZN (n_0), .A1 (n_34), .A2 (p_1[30]), .B1 (p_0[30]), .B2 (n_33));
XNOR2_X1 i_0 (.ZN (p_2[30]), .A (n_32), .B (n_0));
FA_X1 i_29 (.CO (n_29), .S (p_2[28]), .A (p_0[28]), .B (p_1[28]), .CI (n_28));
FA_X1 i_28 (.CO (n_28), .S (p_2[27]), .A (p_0[27]), .B (p_1[27]), .CI (n_27));
FA_X1 i_27 (.CO (n_27), .S (p_2[26]), .A (p_0[26]), .B (p_1[26]), .CI (slo__sro_n269));
INV_X1 slo__sro_c202 (.ZN (slo__sro_n289), .A (n_23));
NOR2_X1 slo__sro_c553 (.ZN (slo__sro_n776), .A1 (p_1[10]), .A2 (p_0[10]));
INV_X1 slo__sro_c216 (.ZN (slo__sro_n306), .A (n_16));
NAND2_X2 slo__sro_c449 (.ZN (slo__sro_n603), .A1 (slo__sro_n286), .A2 (p_1[24]));
FA_X1 i_22 (.CO (n_22), .S (p_2[21]), .A (p_0[21]), .B (p_1[21]), .CI (n_21));
FA_X1 i_21 (.CO (n_21), .S (p_2[20]), .A (p_0[20]), .B (p_1[20]), .CI (n_20));
FA_X1 i_20 (.CO (n_20), .S (p_2[19]), .A (p_0[19]), .B (p_1[19]), .CI (n_19));
FA_X1 i_19 (.CO (n_19), .S (p_2[18]), .A (p_0[18]), .B (p_1[18]), .CI (n_18));
FA_X1 i_18 (.CO (n_18), .S (p_2[17]), .A (p_0[17]), .B (p_1[17]), .CI (slo__sro_n303));
INV_X1 slo__sro_c267 (.ZN (slo__sro_n386), .A (p_1[2]));
FA_X1 i_16 (.CO (n_16), .S (p_2[15]), .A (p_0[15]), .B (p_1[15]), .CI (CLOCK_slo__sro_n1110));
FA_X1 i_14 (.CO (n_14), .S (p_2[13]), .A (p_0[13]), .B (p_1[13]), .CI (n_13));
FA_X1 i_13 (.CO (n_13), .S (p_2[12]), .A (p_0[12]), .B (p_1[12]), .CI (slo__sro_n252));
OAI21_X2 slo__sro_c270 (.ZN (n_3), .A (slo__sro_n385), .B1 (slo__sro_n384), .B2 (slo__sro_n386));
INV_X1 CLOCK_slo__sro_c677 (.ZN (CLOCK_slo__sro_n998), .A (p_0[0]));
FA_X1 i_10 (.CO (n_10), .S (p_2[9]), .A (p_0[9]), .B (p_1[9]), .CI (slo__sro_n164));
INV_X1 slo__sro_c188 (.ZN (slo__sro_n272), .A (slo__sro_n602));
FA_X1 i_8 (.CO (n_8), .S (p_2[7]), .A (p_0[7]), .B (p_1[7]), .CI (n_7));
FA_X1 i_7 (.CO (n_7), .S (p_2[6]), .A (p_0[6]), .B (p_1[6]), .CI (n_6));
FA_X1 i_6 (.CO (n_6), .S (p_2[5]), .A (p_0[5]), .B (p_1[5]), .CI (n_5));
FA_X1 i_5 (.CO (n_5), .S (p_2[4]), .A (p_0[4]), .B (p_1[4]), .CI (n_4));
INV_X2 CLOCK_slo__sro_c796 (.ZN (CLOCK_slo__sro_n1113), .A (n_14));
NAND2_X1 slo__sro_c447 (.ZN (slo__sro_n605), .A1 (p_1[24]), .A2 (p_0[24]));
INV_X2 slo__sro_c95 (.ZN (slo__sro_n167), .A (n_8));
NAND2_X1 CLOCK_slo__sro_c691 (.ZN (CLOCK_slo__sro_n1012), .A1 (p_1[3]), .A2 (p_0[3]));
INV_X1 slo__sro_c42 (.ZN (slo__sro_n111), .A (p_1[1]));
NAND2_X1 slo__sro_c43 (.ZN (slo__sro_n110), .A1 (n_1), .A2 (p_0[1]));
NOR2_X2 slo__sro_c44 (.ZN (slo__sro_n109), .A1 (n_1), .A2 (p_0[1]));
OAI21_X4 slo__sro_c45 (.ZN (slo__sro_n108), .A (slo__sro_n110), .B1 (slo__sro_n109), .B2 (slo__sro_n111));
XNOR2_X1 slo__sro_c46 (.ZN (slo__sro_n107), .A (n_1), .B (p_0[1]));
XNOR2_X1 slo__sro_c47 (.ZN (p_2[1]), .A (slo__sro_n107), .B (p_1[1]));
NAND2_X1 slo__sro_c96 (.ZN (slo__sro_n166), .A1 (p_1[8]), .A2 (p_0[8]));
NOR2_X1 CLOCK_slo__sro_c798 (.ZN (CLOCK_slo__sro_n1111), .A1 (p_1[14]), .A2 (p_0[14]));
OAI21_X2 slo__sro_c98 (.ZN (slo__sro_n164), .A (slo__sro_n166), .B1 (slo__sro_n167), .B2 (CLOCK_slo__mro_n1049));
INV_X1 slo__sro_c551 (.ZN (slo__sro_n778), .A (n_10));
NAND2_X1 slo__sro_c552 (.ZN (slo__sro_n777), .A1 (p_1[10]), .A2 (p_0[10]));
NAND2_X1 slo__sro_c189 (.ZN (slo__sro_n271), .A1 (p_1[25]), .A2 (p_0[25]));
NOR2_X1 slo__sro_c190 (.ZN (slo__sro_n270), .A1 (p_1[25]), .A2 (p_0[25]));
OAI21_X1 slo__sro_c191 (.ZN (slo__sro_n269), .A (slo__sro_n271), .B1 (slo__sro_n272), .B2 (slo__sro_n270));
XNOR2_X2 slo__sro_c192 (.ZN (slo__sro_n268), .A (p_1[25]), .B (p_0[25]));
XNOR2_X2 slo__sro_c193 (.ZN (p_2[25]), .A (slo__sro_n268), .B (slo__sro_n602));
NAND2_X1 slo__sro_c203 (.ZN (slo__sro_n288), .A1 (p_1[23]), .A2 (p_0[23]));
NOR2_X1 slo__sro_c204 (.ZN (slo__sro_n287), .A1 (p_1[23]), .A2 (p_0[23]));
OAI21_X4 slo__sro_c205 (.ZN (slo__sro_n286), .A (slo__sro_n288), .B1 (slo__sro_n289), .B2 (slo__sro_n287));
XNOR2_X1 slo__sro_c206 (.ZN (slo__sro_n285), .A (p_1[23]), .B (p_0[23]));
XNOR2_X2 slo__sro_c207 (.ZN (p_2[23]), .A (slo__sro_n285), .B (n_23));
NAND2_X1 slo__sro_c217 (.ZN (slo__sro_n305), .A1 (p_1[16]), .A2 (p_0[16]));
NOR2_X1 slo__sro_c218 (.ZN (slo__sro_n304), .A1 (p_1[16]), .A2 (p_0[16]));
OAI21_X1 slo__sro_c219 (.ZN (slo__sro_n303), .A (slo__sro_n305), .B1 (slo__sro_n304), .B2 (slo__sro_n306));
XNOR2_X1 slo__sro_c220 (.ZN (slo__sro_n302), .A (p_1[16]), .B (p_0[16]));
XNOR2_X1 slo__sro_c221 (.ZN (p_2[16]), .A (slo__sro_n302), .B (n_16));
NAND2_X1 slo__sro_c268 (.ZN (slo__sro_n385), .A1 (slo__sro_n108), .A2 (p_0[2]));
NOR2_X1 slo__sro_c269 (.ZN (slo__sro_n384), .A1 (slo__sro_n108), .A2 (p_0[2]));
INV_X1 slo__sro_c174 (.ZN (slo__sro_n255), .A (slo__sro_n775));
NAND2_X1 slo__sro_c175 (.ZN (slo__sro_n254), .A1 (p_1[11]), .A2 (p_0[11]));
NOR2_X1 slo__sro_c176 (.ZN (slo__sro_n253), .A1 (p_1[11]), .A2 (p_0[11]));
OAI21_X1 slo__sro_c177 (.ZN (slo__sro_n252), .A (slo__sro_n254), .B1 (slo__sro_n255), .B2 (slo__sro_n253));
XNOR2_X1 slo__sro_c178 (.ZN (slo__sro_n251), .A (p_1[11]), .B (p_0[11]));
XNOR2_X1 slo__sro_c179 (.ZN (p_2[11]), .A (slo__sro_n251), .B (slo__sro_n775));
XNOR2_X2 slo__sro_c271 (.ZN (slo__sro_n383), .A (slo__sro_n108), .B (p_0[2]));
XNOR2_X1 slo__sro_c272 (.ZN (p_2[2]), .A (slo__sro_n383), .B (p_1[2]));
NAND2_X2 slo__sro_c448 (.ZN (slo__sro_n604), .A1 (slo__sro_n286), .A2 (p_0[24]));
INV_X1 slo__sro_c306 (.ZN (slo__sro_n426), .A (n_22));
NAND2_X1 slo__sro_c307 (.ZN (slo__sro_n425), .A1 (p_1[22]), .A2 (p_0[22]));
NOR2_X1 slo__sro_c308 (.ZN (slo__sro_n424), .A1 (p_1[22]), .A2 (p_0[22]));
OAI21_X2 slo__sro_c309 (.ZN (n_23), .A (slo__sro_n425), .B1 (slo__sro_n426), .B2 (slo__sro_n424));
XNOR2_X1 slo__sro_c310 (.ZN (slo__sro_n423), .A (p_1[22]), .B (p_0[22]));
XNOR2_X1 slo__sro_c311 (.ZN (p_2[22]), .A (slo__sro_n423), .B (n_22));
NAND3_X4 slo__sro_c450 (.ZN (slo__sro_n602), .A1 (slo__sro_n604), .A2 (slo__sro_n603), .A3 (slo__sro_n605));
XNOR2_X1 slo__sro_c451 (.ZN (slo__sro_n601), .A (p_1[24]), .B (p_0[24]));
XNOR2_X1 slo__sro_c452 (.ZN (p_2[24]), .A (slo__sro_n601), .B (slo__sro_n286));
OAI21_X1 slo__sro_c554 (.ZN (slo__sro_n775), .A (slo__sro_n777), .B1 (slo__sro_n778), .B2 (slo__sro_n776));
XNOR2_X1 slo__sro_c555 (.ZN (slo__sro_n774), .A (p_1[10]), .B (p_0[10]));
XNOR2_X1 slo__sro_c556 (.ZN (p_2[10]), .A (slo__sro_n774), .B (n_10));
XNOR2_X1 slo__mro_c541 (.ZN (slo__mro_n761), .A (p_1[8]), .B (p_0[8]));
XNOR2_X1 slo__mro_c542 (.ZN (p_2[8]), .A (n_8), .B (slo__mro_n761));
INV_X1 slo__sro_c514 (.ZN (slo__sro_n726), .A (n_30));
NOR2_X1 slo__sro_c515 (.ZN (slo__sro_n725), .A1 (n_33), .A2 (p_0[30]));
NAND2_X1 slo__sro_c516 (.ZN (slo__sro_n724), .A1 (slo__sro_n725), .A2 (slo__sro_n726));
OR2_X1 slo__sro_c517 (.ZN (slo__sro_n723), .A1 (p_1[30]), .A2 (n_34));
OAI21_X1 slo__sro_c518 (.ZN (n_31), .A (slo__sro_n724), .B1 (n_32), .B2 (slo__sro_n723));
NOR2_X2 CLOCK_slo__sro_c679 (.ZN (n_1), .A1 (CLOCK_slo__sro_n997), .A2 (CLOCK_slo__sro_n998));
XNOR2_X1 CLOCK_slo__sro_c680 (.ZN (p_2[0]), .A (p_1[0]), .B (CLOCK_slo__sro_n998));
OAI21_X1 CLOCK_slo__sro_c692 (.ZN (CLOCK_slo__sro_n1011), .A (n_3), .B1 (p_1[3]), .B2 (p_0[3]));
NAND2_X1 CLOCK_slo__sro_c693 (.ZN (n_4), .A1 (CLOCK_slo__sro_n1012), .A2 (CLOCK_slo__sro_n1011));
XNOR2_X2 CLOCK_slo__sro_c694 (.ZN (CLOCK_slo__sro_n1010), .A (p_1[3]), .B (p_0[3]));
XNOR2_X2 CLOCK_slo__sro_c695 (.ZN (p_2[3]), .A (CLOCK_slo__sro_n1010), .B (n_3));
NAND2_X1 CLOCK_slo__sro_c797 (.ZN (CLOCK_slo__sro_n1112), .A1 (p_1[14]), .A2 (p_0[14]));
NOR2_X1 CLOCK_slo__mro_c743 (.ZN (CLOCK_slo__mro_n1049), .A1 (p_1[8]), .A2 (p_0[8]));
OAI21_X2 CLOCK_slo__sro_c799 (.ZN (CLOCK_slo__sro_n1110), .A (CLOCK_slo__sro_n1112)
    , .B1 (CLOCK_slo__sro_n1113), .B2 (CLOCK_slo__sro_n1111));
XNOR2_X1 CLOCK_slo__sro_c800 (.ZN (CLOCK_slo__sro_n1109), .A (p_1[14]), .B (p_0[14]));
XNOR2_X1 CLOCK_slo__sro_c801 (.ZN (p_2[14]), .A (CLOCK_slo__sro_n1109), .B (n_14));
INV_X1 CLOCK_slo__sro_c829 (.ZN (CLOCK_slo__sro_n1148), .A (n_29));
NAND2_X1 CLOCK_slo__sro_c830 (.ZN (CLOCK_slo__sro_n1147), .A1 (p_1[29]), .A2 (p_0[29]));
NOR2_X1 CLOCK_slo__sro_c831 (.ZN (CLOCK_slo__sro_n1146), .A1 (p_1[29]), .A2 (p_0[29]));
OAI21_X1 CLOCK_slo__sro_c832 (.ZN (n_30), .A (CLOCK_slo__sro_n1147), .B1 (CLOCK_slo__sro_n1148), .B2 (CLOCK_slo__sro_n1146));
XNOR2_X1 CLOCK_slo__sro_c833 (.ZN (CLOCK_slo__sro_n1145), .A (p_1[29]), .B (p_0[29]));
XNOR2_X1 CLOCK_slo__sro_c834 (.ZN (p_2[29]), .A (n_29), .B (CLOCK_slo__sro_n1145));

endmodule //datapath__0_127

module datapath__0_126 (Multiplier, p_0, p_1);

output [31:0] p_1;
input [31:0] Multiplier;
input [31:0] p_0;
wire slo__sro_n770;
wire slo__sro_n740;
wire n_1;
wire n_2;
wire n_3;
wire slo__sro_n406;
wire n_5;
wire n_6;
wire n_8;
wire n_9;
wire n_10;
wire n_12;
wire n_13;
wire n_14;
wire n_15;
wire n_16;
wire n_17;
wire n_19;
wire n_20;
wire n_21;
wire CLOCK_slo__sro_n985;
wire n_23;
wire n_25;
wire n_26;
wire n_27;
wire n_28;
wire n_29;
wire n_30;
wire n_32;
wire n_0;
wire n_34;
wire n_33;
wire n_31;
wire slo__sro_n99;
wire slo__sro_n100;
wire slo__sro_n101;
wire slo__sro_n102;
wire slo__sro_n103;
wire slo__sro_n116;
wire slo__sro_n117;
wire slo__sro_n118;
wire slo__sro_n119;
wire slo__sro_n402;
wire slo__sro_n403;
wire slo__sro_n404;
wire slo__sro_n405;
wire slo__sro_n144;
wire slo__sro_n145;
wire slo__sro_n146;
wire slo__sro_n147;
wire slo__sro_n148;
wire slo__sro_n546;
wire slo__sro_n547;
wire slo__sro_n548;
wire slo__sro_n549;
wire slo__sro_n741;
wire slo__sro_n742;
wire slo__sro_n743;
wire CLOCK_slo__sro_n1053;
wire slo__sro_n612;
wire slo__sro_n613;
wire slo__sro_n614;
wire slo__sro_n771;
wire slo__sro_n772;
wire slo__sro_n773;
wire slo__sro_n774;
wire CLOCK_slo__sro_n954;
wire CLOCK_slo__sro_n955;
wire CLOCK_slo__sro_n956;
wire CLOCK_slo__sro_n957;
wire slo__sro_n275;
wire slo__sro_n276;
wire slo__sro_n277;
wire slo__sro_n278;
wire slo__sro_n279;
wire CLOCK_slo__sro_n986;
wire CLOCK_slo__sro_n987;
wire CLOCK_slo__sro_n988;
wire CLOCK_slo__sro_n1006;
wire CLOCK_slo__sro_n1007;
wire CLOCK_slo__sro_n1008;
wire CLOCK_slo__sro_n1009;
wire CLOCK_slo__sro_n1010;
wire CLOCK_slo__mro_n1023;
wire CLOCK_slo__sro_n1054;
wire CLOCK_slo__sro_n1055;
wire CLOCK_slo__sro_n1056;


INV_X1 i_36 (.ZN (n_34), .A (Multiplier[30]));
INV_X1 i_35 (.ZN (n_33), .A (p_0[30]));
INV_X1 i_34 (.ZN (n_32), .A (n_30));
OAI33_X1 i_33 (.ZN (n_31), .A1 (n_32), .A2 (p_0[30]), .A3 (n_34), .B1 (n_30), .B2 (n_33), .B3 (Multiplier[30]));
XOR2_X1 i_32 (.Z (p_1[31]), .A (Multiplier[31]), .B (n_31));
OAI22_X1 i_31 (.ZN (n_0), .A1 (n_34), .A2 (p_0[30]), .B1 (Multiplier[30]), .B2 (n_33));
XNOR2_X1 i_0 (.ZN (p_1[30]), .A (n_32), .B (n_0));
FA_X1 i_30 (.CO (n_30), .S (p_1[29]), .A (Multiplier[29]), .B (p_0[29]), .CI (n_29));
NAND2_X1 slo__sro_c592 (.ZN (slo__sro_n773), .A1 (p_0[10]), .A2 (Multiplier[10]));
INV_X2 slo__sro_c591 (.ZN (slo__sro_n774), .A (n_10));
INV_X1 slo__sro_c564 (.ZN (slo__sro_n743), .A (n_27));
FA_X1 i_26 (.CO (n_26), .S (p_1[25]), .A (Multiplier[25]), .B (p_0[25]), .CI (n_25));
FA_X1 i_25 (.CO (n_25), .S (p_1[24]), .A (Multiplier[24]), .B (p_0[24]), .CI (slo__sro_n100));
INV_X1 slo__sro_c54 (.ZN (slo__sro_n119), .A (n_26));
NOR2_X1 slo__sro_c566 (.ZN (slo__sro_n741), .A1 (p_0[27]), .A2 (Multiplier[27]));
XNOR2_X1 CLOCK_slo__sro_c691 (.ZN (p_1[2]), .A (CLOCK_slo__sro_n954), .B (n_2));
INV_X1 CLOCK_slo__sro_c737 (.ZN (CLOCK_slo__sro_n1010), .A (n_17));
FA_X1 i_20 (.CO (n_20), .S (p_1[19]), .A (Multiplier[19]), .B (p_0[19]), .CI (n_19));
FA_X1 i_19 (.CO (n_19), .S (p_1[18]), .A (Multiplier[18]), .B (p_0[18]), .CI (CLOCK_slo__sro_n1007));
XNOR2_X1 CLOCK_slo__mro_c751 (.ZN (CLOCK_slo__mro_n1023), .A (n_28), .B (Multiplier[28]));
FA_X1 i_17 (.CO (n_17), .S (p_1[16]), .A (Multiplier[16]), .B (p_0[16]), .CI (n_16));
FA_X1 i_16 (.CO (n_16), .S (p_1[15]), .A (Multiplier[15]), .B (p_0[15]), .CI (n_15));
FA_X1 i_15 (.CO (n_15), .S (p_1[14]), .A (Multiplier[14]), .B (p_0[14]), .CI (n_14));
FA_X1 i_14 (.CO (n_14), .S (p_1[13]), .A (Multiplier[13]), .B (p_0[13]), .CI (n_13));
FA_X1 i_13 (.CO (n_13), .S (p_1[12]), .A (Multiplier[12]), .B (p_0[12]), .CI (n_12));
INV_X1 CLOCK_slo__sro_c686 (.ZN (CLOCK_slo__sro_n957), .A (n_2));
FA_X1 i_10 (.CO (n_10), .S (p_1[9]), .A (Multiplier[9]), .B (p_0[9]), .CI (n_9));
FA_X1 i_9 (.CO (n_9), .S (p_1[8]), .A (Multiplier[8]), .B (p_0[8]), .CI (n_8));
FA_X1 i_8 (.CO (n_8), .S (p_1[7]), .A (Multiplier[7]), .B (p_0[7]), .CI (slo__sro_n403));
NAND2_X1 slo__sro_c565 (.ZN (slo__sro_n742), .A1 (p_0[27]), .A2 (Multiplier[27]));
FA_X1 i_6 (.CO (n_6), .S (p_1[5]), .A (Multiplier[5]), .B (p_0[5]), .CI (n_5));
FA_X1 i_5 (.CO (n_5), .S (p_1[4]), .A (Multiplier[4]), .B (p_0[4]), .CI (slo__sro_n145));
XNOR2_X2 slo__sro_c303 (.ZN (p_1[6]), .A (slo__sro_n402), .B (n_6));
INV_X1 CLOCK_slo__sro_c717 (.ZN (CLOCK_slo__sro_n988), .A (n_20));
FA_X1 i_2 (.CO (n_2), .S (p_1[1]), .A (Multiplier[1]), .B (p_0[1]), .CI (n_1));
HA_X1 i_1 (.CO (n_1), .S (p_1[0]), .A (Multiplier[0]), .B (p_0[0]));
INV_X1 slo__sro_c40 (.ZN (slo__sro_n103), .A (n_23));
NAND2_X1 slo__sro_c41 (.ZN (slo__sro_n102), .A1 (p_0[23]), .A2 (Multiplier[23]));
NOR2_X1 slo__sro_c42 (.ZN (slo__sro_n101), .A1 (p_0[23]), .A2 (Multiplier[23]));
OAI21_X1 slo__sro_c43 (.ZN (slo__sro_n100), .A (slo__sro_n102), .B1 (slo__sro_n103), .B2 (slo__sro_n101));
XNOR2_X2 slo__sro_c44 (.ZN (slo__sro_n99), .A (p_0[23]), .B (Multiplier[23]));
XNOR2_X2 slo__sro_c45 (.ZN (p_1[23]), .A (slo__sro_n99), .B (n_23));
NAND2_X1 slo__sro_c55 (.ZN (slo__sro_n118), .A1 (p_0[26]), .A2 (Multiplier[26]));
NOR2_X1 slo__sro_c56 (.ZN (slo__sro_n117), .A1 (p_0[26]), .A2 (Multiplier[26]));
OAI21_X2 slo__sro_c57 (.ZN (n_27), .A (slo__sro_n118), .B1 (slo__sro_n119), .B2 (slo__sro_n117));
XNOR2_X1 slo__sro_c58 (.ZN (slo__sro_n116), .A (p_0[26]), .B (Multiplier[26]));
XNOR2_X1 slo__sro_c59 (.ZN (p_1[26]), .A (n_26), .B (slo__sro_n116));
INV_X1 slo__sro_c298 (.ZN (slo__sro_n406), .A (n_6));
NAND2_X1 slo__sro_c299 (.ZN (slo__sro_n405), .A1 (p_0[6]), .A2 (Multiplier[6]));
NOR2_X1 slo__sro_c300 (.ZN (slo__sro_n404), .A1 (p_0[6]), .A2 (Multiplier[6]));
OAI21_X2 slo__sro_c301 (.ZN (slo__sro_n403), .A (slo__sro_n405), .B1 (slo__sro_n406), .B2 (slo__sro_n404));
XNOR2_X2 slo__sro_c302 (.ZN (slo__sro_n402), .A (p_0[6]), .B (Multiplier[6]));
INV_X1 slo__sro_c81 (.ZN (slo__sro_n148), .A (n_3));
NAND2_X1 slo__sro_c82 (.ZN (slo__sro_n147), .A1 (p_0[3]), .A2 (Multiplier[3]));
NOR2_X1 slo__sro_c83 (.ZN (slo__sro_n146), .A1 (p_0[3]), .A2 (Multiplier[3]));
OAI21_X1 slo__sro_c84 (.ZN (slo__sro_n145), .A (slo__sro_n147), .B1 (slo__sro_n148), .B2 (slo__sro_n146));
XNOR2_X1 slo__sro_c85 (.ZN (slo__sro_n144), .A (p_0[3]), .B (Multiplier[3]));
XNOR2_X1 slo__sro_c86 (.ZN (p_1[3]), .A (n_3), .B (slo__sro_n144));
INV_X1 slo__sro_c410 (.ZN (slo__sro_n549), .A (slo__sro_n276));
NAND2_X1 slo__sro_c411 (.ZN (slo__sro_n548), .A1 (p_0[22]), .A2 (Multiplier[22]));
NOR2_X1 slo__sro_c412 (.ZN (slo__sro_n547), .A1 (p_0[22]), .A2 (Multiplier[22]));
OAI21_X2 slo__sro_c413 (.ZN (n_23), .A (slo__sro_n548), .B1 (slo__sro_n549), .B2 (slo__sro_n547));
XNOR2_X2 slo__sro_c414 (.ZN (slo__sro_n546), .A (p_0[22]), .B (Multiplier[22]));
XNOR2_X2 slo__sro_c415 (.ZN (p_1[22]), .A (slo__sro_n546), .B (slo__sro_n276));
OAI21_X2 slo__sro_c567 (.ZN (n_28), .A (slo__sro_n742), .B1 (slo__sro_n743), .B2 (slo__sro_n741));
XNOR2_X2 slo__sro_c568 (.ZN (slo__sro_n740), .A (p_0[27]), .B (Multiplier[27]));
XNOR2_X1 slo__sro_c569 (.ZN (p_1[27]), .A (n_27), .B (slo__sro_n740));
INV_X1 slo__sro_c471 (.ZN (slo__sro_n614), .A (n_28));
NAND2_X1 slo__sro_c472 (.ZN (slo__sro_n613), .A1 (p_0[28]), .A2 (Multiplier[28]));
NOR2_X1 slo__sro_c473 (.ZN (slo__sro_n612), .A1 (p_0[28]), .A2 (Multiplier[28]));
OAI21_X1 slo__sro_c474 (.ZN (n_29), .A (slo__sro_n613), .B1 (slo__sro_n612), .B2 (slo__sro_n614));
INV_X1 CLOCK_slo__sro_c779 (.ZN (CLOCK_slo__sro_n1056), .A (slo__sro_n771));
NAND2_X1 CLOCK_slo__sro_c780 (.ZN (CLOCK_slo__sro_n1055), .A1 (p_0[11]), .A2 (Multiplier[11]));
NOR2_X1 slo__sro_c593 (.ZN (slo__sro_n772), .A1 (p_0[10]), .A2 (Multiplier[10]));
OAI21_X2 slo__sro_c594 (.ZN (slo__sro_n771), .A (slo__sro_n773), .B1 (slo__sro_n774), .B2 (slo__sro_n772));
XNOR2_X1 slo__sro_c595 (.ZN (slo__sro_n770), .A (p_0[10]), .B (Multiplier[10]));
XNOR2_X1 slo__sro_c596 (.ZN (p_1[10]), .A (slo__sro_n770), .B (n_10));
NAND2_X1 CLOCK_slo__sro_c687 (.ZN (CLOCK_slo__sro_n956), .A1 (p_0[2]), .A2 (Multiplier[2]));
NOR2_X1 CLOCK_slo__sro_c688 (.ZN (CLOCK_slo__sro_n955), .A1 (p_0[2]), .A2 (Multiplier[2]));
OAI21_X1 CLOCK_slo__sro_c689 (.ZN (n_3), .A (CLOCK_slo__sro_n956), .B1 (CLOCK_slo__sro_n957), .B2 (CLOCK_slo__sro_n955));
XNOR2_X1 CLOCK_slo__sro_c690 (.ZN (CLOCK_slo__sro_n954), .A (p_0[2]), .B (Multiplier[2]));
INV_X2 slo__sro_c199 (.ZN (slo__sro_n279), .A (n_21));
NAND2_X1 slo__sro_c200 (.ZN (slo__sro_n278), .A1 (p_0[21]), .A2 (Multiplier[21]));
NOR2_X1 slo__sro_c201 (.ZN (slo__sro_n277), .A1 (p_0[21]), .A2 (Multiplier[21]));
OAI21_X2 slo__sro_c202 (.ZN (slo__sro_n276), .A (slo__sro_n278), .B1 (slo__sro_n279), .B2 (slo__sro_n277));
XNOR2_X2 slo__sro_c203 (.ZN (slo__sro_n275), .A (p_0[21]), .B (Multiplier[21]));
XNOR2_X2 slo__sro_c204 (.ZN (p_1[21]), .A (n_21), .B (slo__sro_n275));
NAND2_X1 CLOCK_slo__sro_c718 (.ZN (CLOCK_slo__sro_n987), .A1 (p_0[20]), .A2 (Multiplier[20]));
NOR2_X1 CLOCK_slo__sro_c719 (.ZN (CLOCK_slo__sro_n986), .A1 (p_0[20]), .A2 (Multiplier[20]));
OAI21_X1 CLOCK_slo__sro_c720 (.ZN (n_21), .A (CLOCK_slo__sro_n987), .B1 (CLOCK_slo__sro_n988), .B2 (CLOCK_slo__sro_n986));
XNOR2_X1 CLOCK_slo__sro_c721 (.ZN (CLOCK_slo__sro_n985), .A (p_0[20]), .B (Multiplier[20]));
XNOR2_X1 CLOCK_slo__sro_c722 (.ZN (p_1[20]), .A (n_20), .B (CLOCK_slo__sro_n985));
NAND2_X1 CLOCK_slo__sro_c738 (.ZN (CLOCK_slo__sro_n1009), .A1 (p_0[17]), .A2 (Multiplier[17]));
NOR2_X1 CLOCK_slo__sro_c739 (.ZN (CLOCK_slo__sro_n1008), .A1 (p_0[17]), .A2 (Multiplier[17]));
OAI21_X1 CLOCK_slo__sro_c740 (.ZN (CLOCK_slo__sro_n1007), .A (CLOCK_slo__sro_n1009)
    , .B1 (CLOCK_slo__sro_n1010), .B2 (CLOCK_slo__sro_n1008));
XNOR2_X1 CLOCK_slo__sro_c741 (.ZN (CLOCK_slo__sro_n1006), .A (p_0[17]), .B (Multiplier[17]));
XNOR2_X1 CLOCK_slo__sro_c742 (.ZN (p_1[17]), .A (n_17), .B (CLOCK_slo__sro_n1006));
XNOR2_X1 CLOCK_slo__mro_c752 (.ZN (p_1[28]), .A (CLOCK_slo__mro_n1023), .B (p_0[28]));
NOR2_X1 CLOCK_slo__sro_c781 (.ZN (CLOCK_slo__sro_n1054), .A1 (p_0[11]), .A2 (Multiplier[11]));
OAI21_X1 CLOCK_slo__sro_c782 (.ZN (n_12), .A (CLOCK_slo__sro_n1055), .B1 (CLOCK_slo__sro_n1056), .B2 (CLOCK_slo__sro_n1054));
XNOR2_X1 CLOCK_slo__sro_c783 (.ZN (CLOCK_slo__sro_n1053), .A (p_0[11]), .B (Multiplier[11]));
XNOR2_X1 CLOCK_slo__sro_c784 (.ZN (p_1[11]), .A (CLOCK_slo__sro_n1053), .B (slo__sro_n771));

endmodule //datapath__0_126

module datapath__0_122 (p_0, p_1, p_2);

output [31:0] p_2;
input [31:0] p_0;
input [31:0] p_1;
wire CLOCK_slo__sro_n1166;
wire slo__sro_n464;
wire CLOCK_slo__mro_n1149;
wire slo__sro_n669;
wire n_1;
wire n_2;
wire slo__sro_n319;
wire n_8;
wire n_9;
wire n_10;
wire n_11;
wire n_14;
wire n_15;
wire n_18;
wire n_19;
wire n_20;
wire n_21;
wire n_22;
wire n_23;
wire n_24;
wire n_27;
wire n_29;
wire n_30;
wire n_32;
wire n_0;
wire n_34;
wire n_33;
wire n_31;
wire slo__sro_n138;
wire slo__sro_n139;
wire slo__sro_n140;
wire slo__sro_n141;
wire slo__sro_n142;
wire slo__n893;
wire slo__sro_n156;
wire slo__sro_n157;
wire slo__sro_n158;
wire slo__sro_n159;
wire slo__sro_n189;
wire slo__sro_n190;
wire slo__sro_n191;
wire slo__sro_n192;
wire slo__sro_n202;
wire slo__sro_n203;
wire slo__sro_n204;
wire slo__sro_n205;
wire slo__sro_n217;
wire slo__sro_n218;
wire slo__sro_n219;
wire slo__sro_n220;
wire slo__sro_n221;
wire slo__sro_n273;
wire slo__sro_n274;
wire slo__sro_n275;
wire slo__sro_n276;
wire slo__sro_n277;
wire slo__sro_n320;
wire slo__sro_n321;
wire slo__sro_n322;
wire slo__sro_n365;
wire slo__sro_n366;
wire slo__sro_n367;
wire slo__sro_n368;
wire slo__sro_n407;
wire slo__sro_n408;
wire slo__sro_n409;
wire slo__sro_n410;
wire slo__sro_n411;
wire slo__sro_n465;
wire slo__sro_n466;
wire slo__sro_n467;
wire slo__sro_n468;
wire slo__sro_n636;
wire slo__sro_n637;
wire slo__sro_n638;
wire slo__sro_n639;
wire slo__sro_n498;
wire slo__sro_n499;
wire slo__sro_n500;
wire slo__sro_n501;
wire slo__sro_n670;
wire slo__sro_n671;
wire slo__sro_n672;
wire slo__sro_n712;
wire slo__sro_n713;
wire slo__sro_n714;
wire slo__sro_n715;
wire slo__sro_n716;
wire slo__sro_n733;
wire slo__sro_n734;
wire slo__sro_n735;
wire slo__sro_n736;
wire slo__sro_n737;
wire slo__mro_n765;
wire CLOCK_slo__mro_n1112;
wire CLOCK_slo__sro_n1167;
wire CLOCK_slo__sro_n1168;
wire CLOCK_slo__sro_n1169;
wire CLOCK_slo__sro_n1195;
wire CLOCK_slo__sro_n1196;
wire CLOCK_slo__sro_n1197;
wire CLOCK_slo__sro_n1198;
wire CLOCK_slo__sro_n1199;


INV_X1 i_36 (.ZN (n_34), .A (p_0[30]));
INV_X1 i_35 (.ZN (n_33), .A (p_1[30]));
INV_X1 i_34 (.ZN (n_32), .A (n_30));
OAI33_X1 i_33 (.ZN (n_31), .A1 (n_34), .A2 (p_1[30]), .A3 (n_32), .B1 (n_30), .B2 (n_33), .B3 (p_0[30]));
XOR2_X1 i_32 (.Z (p_2[31]), .A (p_0[31]), .B (n_31));
OAI22_X1 i_31 (.ZN (n_0), .A1 (n_34), .A2 (p_1[30]), .B1 (p_0[30]), .B2 (n_33));
XNOR2_X1 i_0 (.ZN (p_2[30]), .A (n_32), .B (n_0));
FA_X1 i_30 (.CO (n_30), .S (p_2[29]), .A (p_0[29]), .B (p_1[29]), .CI (n_29));
INV_X2 slo__sro_c137 (.ZN (slo__sro_n221), .A (n_15));
INV_X1 slo__sro_c255 (.ZN (slo__sro_n411), .A (CLOCK_slo__sro_n1196));
INV_X1 slo__sro_c229 (.ZN (slo__sro_n368), .A (p_1[27]));
NAND2_X1 slo__sro_c301 (.ZN (slo__sro_n467), .A1 (p_1[12]), .A2 (p_0[12]));
FA_X1 i_24 (.CO (n_24), .S (p_2[23]), .A (p_0[23]), .B (p_1[23]), .CI (n_23));
FA_X1 i_23 (.CO (n_23), .S (p_2[22]), .A (p_0[22]), .B (p_1[22]), .CI (n_22));
FA_X1 i_22 (.CO (n_22), .S (p_2[21]), .A (p_0[21]), .B (p_1[21]), .CI (n_21));
INV_X1 slo__sro_c123 (.ZN (slo__sro_n205), .A (slo__sro_n365));
FA_X1 i_20 (.CO (n_20), .S (p_2[19]), .A (p_0[19]), .B (p_1[19]), .CI (n_19));
FA_X1 i_19 (.CO (n_19), .S (p_2[18]), .A (p_0[18]), .B (p_1[18]), .CI (n_18));
FA_X1 i_18 (.CO (n_18), .S (p_2[17]), .A (p_0[17]), .B (p_1[17]), .CI (slo__sro_n637));
NAND2_X1 slo__sro_c445 (.ZN (slo__sro_n672), .A1 (p_1[4]), .A2 (p_0[4]));
INV_X1 slo__sro_c300 (.ZN (slo__sro_n468), .A (slo__sro_n713));
FA_X1 i_15 (.CO (n_15), .S (p_2[14]), .A (p_0[14]), .B (p_1[14]), .CI (n_14));
FA_X1 i_14 (.CO (n_14), .S (p_2[13]), .A (p_0[13]), .B (p_1[13]), .CI (slo__sro_n465));
NAND2_X1 slo__sro_c418 (.ZN (slo__sro_n639), .A1 (slo__sro_n218), .A2 (p_0[16]));
NAND2_X1 slo__sro_c490 (.ZN (slo__sro_n737), .A1 (p_1[5]), .A2 (p_0[5]));
NAND2_X1 slo__sro_c447 (.ZN (slo__sro_n670), .A1 (p_1[4]), .A2 (slo__sro_n139));
FA_X1 i_10 (.CO (n_10), .S (p_2[9]), .A (p_0[9]), .B (p_1[9]), .CI (n_9));
FA_X1 i_8 (.CO (n_8), .S (p_2[7]), .A (p_0[7]), .B (p_1[7]), .CI (slo__sro_n156));
INV_X1 slo__sro_c109 (.ZN (slo__sro_n192), .A (n_20));
XNOR2_X1 slo__mro_c517 (.ZN (slo__mro_n765), .A (slo__sro_n734), .B (p_0[6]));
NAND2_X1 slo__sro_c474 (.ZN (slo__sro_n716), .A1 (p_1[11]), .A2 (p_0[11]));
INV_X1 slo__sro_c80 (.ZN (slo__sro_n159), .A (slo__sro_n734));
NAND2_X1 slo__sro_c208 (.ZN (slo__sro_n321), .A1 (p_1[26]), .A2 (p_0[26]));
FA_X1 i_2 (.CO (n_2), .S (p_2[1]), .A (p_0[1]), .B (p_1[1]), .CI (n_1));
HA_X1 i_1 (.CO (n_1), .S (p_2[0]), .A (p_0[0]), .B (p_1[0]));
INV_X2 slo__sro_c66 (.ZN (slo__sro_n142), .A (slo__sro_n274));
NAND2_X1 slo__sro_c67 (.ZN (slo__sro_n141), .A1 (p_1[3]), .A2 (p_0[3]));
NOR2_X2 slo__sro_c68 (.ZN (slo__sro_n140), .A1 (p_1[3]), .A2 (p_0[3]));
OAI21_X2 slo__sro_c69 (.ZN (slo__sro_n139), .A (slo__sro_n141), .B1 (slo__sro_n140), .B2 (slo__sro_n142));
XNOR2_X1 slo__sro_c70 (.ZN (slo__sro_n138), .A (p_1[3]), .B (p_0[3]));
XNOR2_X1 slo__sro_c71 (.ZN (p_2[3]), .A (slo__sro_n138), .B (slo__sro_n274));
NAND2_X1 slo__sro_c81 (.ZN (slo__sro_n158), .A1 (p_1[6]), .A2 (p_0[6]));
NOR2_X1 slo__sro_c82 (.ZN (slo__sro_n157), .A1 (p_1[6]), .A2 (p_0[6]));
OAI21_X1 slo__sro_c83 (.ZN (slo__sro_n156), .A (slo__sro_n158), .B1 (slo__sro_n157), .B2 (slo__sro_n159));
OAI21_X1 slo__c580 (.ZN (slo__n893), .A (slo__sro_n410), .B1 (slo__sro_n411), .B2 (slo__sro_n409));
XNOR2_X2 CLOCK_slo__mro_c680 (.ZN (CLOCK_slo__mro_n1112), .A (slo__sro_n139), .B (p_0[4]));
NAND2_X1 slo__sro_c110 (.ZN (slo__sro_n191), .A1 (p_1[20]), .A2 (p_0[20]));
NOR2_X1 slo__sro_c111 (.ZN (slo__sro_n190), .A1 (p_1[20]), .A2 (p_0[20]));
OAI21_X1 slo__sro_c112 (.ZN (n_21), .A (slo__sro_n191), .B1 (slo__sro_n192), .B2 (slo__sro_n190));
XNOR2_X1 slo__sro_c113 (.ZN (slo__sro_n189), .A (p_1[20]), .B (p_0[20]));
XNOR2_X1 slo__sro_c114 (.ZN (p_2[20]), .A (slo__sro_n189), .B (n_20));
NAND2_X1 slo__sro_c124 (.ZN (slo__sro_n204), .A1 (p_1[28]), .A2 (p_0[28]));
NOR2_X1 slo__sro_c125 (.ZN (slo__sro_n203), .A1 (p_1[28]), .A2 (p_0[28]));
OAI21_X1 slo__sro_c126 (.ZN (n_29), .A (slo__sro_n204), .B1 (slo__sro_n205), .B2 (slo__sro_n203));
XNOR2_X1 slo__sro_c127 (.ZN (slo__sro_n202), .A (p_1[28]), .B (p_0[28]));
XNOR2_X1 slo__sro_c128 (.ZN (p_2[28]), .A (slo__sro_n202), .B (slo__sro_n365));
NAND2_X1 slo__sro_c138 (.ZN (slo__sro_n220), .A1 (p_1[15]), .A2 (p_0[15]));
NOR2_X1 slo__sro_c139 (.ZN (slo__sro_n219), .A1 (p_1[15]), .A2 (p_0[15]));
OAI21_X2 slo__sro_c140 (.ZN (slo__sro_n218), .A (slo__sro_n220), .B1 (slo__sro_n221), .B2 (slo__sro_n219));
XNOR2_X1 slo__sro_c141 (.ZN (slo__sro_n217), .A (p_1[15]), .B (p_0[15]));
XNOR2_X1 slo__sro_c142 (.ZN (p_2[15]), .A (slo__sro_n217), .B (n_15));
INV_X1 slo__sro_c207 (.ZN (slo__sro_n322), .A (slo__n893));
INV_X1 slo__sro_c185 (.ZN (slo__sro_n277), .A (n_2));
NAND2_X1 slo__sro_c186 (.ZN (slo__sro_n276), .A1 (p_1[2]), .A2 (p_0[2]));
NOR2_X1 slo__sro_c187 (.ZN (slo__sro_n275), .A1 (p_1[2]), .A2 (p_0[2]));
OAI21_X2 slo__sro_c188 (.ZN (slo__sro_n274), .A (slo__sro_n276), .B1 (slo__sro_n277), .B2 (slo__sro_n275));
XNOR2_X1 slo__sro_c189 (.ZN (slo__sro_n273), .A (p_1[2]), .B (p_0[2]));
XNOR2_X1 slo__sro_c190 (.ZN (p_2[2]), .A (slo__sro_n273), .B (n_2));
NOR2_X2 slo__sro_c209 (.ZN (slo__sro_n320), .A1 (p_1[26]), .A2 (p_0[26]));
OAI21_X2 slo__sro_c210 (.ZN (n_27), .A (slo__sro_n321), .B1 (slo__sro_n320), .B2 (slo__sro_n322));
XNOR2_X1 slo__sro_c211 (.ZN (slo__sro_n319), .A (p_1[26]), .B (p_0[26]));
XNOR2_X1 slo__sro_c212 (.ZN (p_2[26]), .A (slo__sro_n319), .B (slo__sro_n408));
NAND2_X1 slo__sro_c230 (.ZN (slo__sro_n367), .A1 (n_27), .A2 (p_0[27]));
NOR2_X1 slo__sro_c231 (.ZN (slo__sro_n366), .A1 (n_27), .A2 (p_0[27]));
OAI21_X2 slo__sro_c232 (.ZN (slo__sro_n365), .A (slo__sro_n367), .B1 (slo__sro_n368), .B2 (slo__sro_n366));
INV_X1 CLOCK_slo__sro_c738 (.ZN (CLOCK_slo__sro_n1169), .A (n_8));
NAND2_X1 CLOCK_slo__sro_c739 (.ZN (CLOCK_slo__sro_n1168), .A1 (p_1[8]), .A2 (p_0[8]));
NAND2_X1 slo__sro_c256 (.ZN (slo__sro_n410), .A1 (p_1[25]), .A2 (p_0[25]));
NOR2_X1 slo__sro_c257 (.ZN (slo__sro_n409), .A1 (p_1[25]), .A2 (p_0[25]));
OAI21_X1 slo__sro_c258 (.ZN (slo__sro_n408), .A (slo__sro_n410), .B1 (slo__sro_n411), .B2 (slo__sro_n409));
XNOR2_X1 slo__sro_c259 (.ZN (slo__sro_n407), .A (p_1[25]), .B (p_0[25]));
XNOR2_X1 slo__sro_c260 (.ZN (p_2[25]), .A (slo__sro_n407), .B (CLOCK_slo__sro_n1196));
NOR2_X2 slo__sro_c302 (.ZN (slo__sro_n466), .A1 (p_1[12]), .A2 (p_0[12]));
OAI21_X1 slo__sro_c303 (.ZN (slo__sro_n465), .A (slo__sro_n467), .B1 (slo__sro_n466), .B2 (slo__sro_n468));
XNOR2_X1 slo__sro_c304 (.ZN (slo__sro_n464), .A (p_1[12]), .B (p_0[12]));
XNOR2_X1 slo__sro_c305 (.ZN (p_2[12]), .A (slo__sro_n464), .B (slo__sro_n713));
OAI21_X2 slo__sro_c419 (.ZN (slo__sro_n638), .A (p_1[16]), .B1 (slo__sro_n218), .B2 (p_0[16]));
NAND2_X2 slo__sro_c420 (.ZN (slo__sro_n637), .A1 (slo__sro_n638), .A2 (slo__sro_n639));
XNOR2_X1 slo__sro_c421 (.ZN (slo__sro_n636), .A (slo__sro_n218), .B (p_0[16]));
XNOR2_X1 slo__sro_c422 (.ZN (p_2[16]), .A (slo__sro_n636), .B (p_1[16]));
NAND2_X1 slo__sro_c446 (.ZN (slo__sro_n671), .A1 (slo__sro_n139), .A2 (p_0[4]));
INV_X1 slo__sro_c329 (.ZN (slo__sro_n501), .A (n_10));
NAND2_X1 slo__sro_c330 (.ZN (slo__sro_n500), .A1 (p_1[10]), .A2 (p_0[10]));
NOR2_X1 slo__sro_c331 (.ZN (slo__sro_n499), .A1 (p_1[10]), .A2 (p_0[10]));
OAI21_X1 slo__sro_c332 (.ZN (n_11), .A (slo__sro_n500), .B1 (slo__sro_n499), .B2 (slo__sro_n501));
XNOR2_X1 slo__sro_c333 (.ZN (slo__sro_n498), .A (p_1[10]), .B (p_0[10]));
XNOR2_X1 slo__sro_c334 (.ZN (p_2[10]), .A (slo__sro_n498), .B (n_10));
NAND3_X2 slo__sro_c448 (.ZN (slo__sro_n669), .A1 (slo__sro_n670), .A2 (slo__sro_n672), .A3 (slo__sro_n671));
XNOR2_X1 CLOCK_slo__mro_c721 (.ZN (CLOCK_slo__mro_n1149), .A (n_27), .B (p_0[27]));
XNOR2_X1 CLOCK_slo__mro_c722 (.ZN (p_2[27]), .A (CLOCK_slo__mro_n1149), .B (p_1[27]));
NAND2_X1 slo__sro_c475 (.ZN (slo__sro_n715), .A1 (n_11), .A2 (p_0[11]));
NAND2_X1 slo__sro_c476 (.ZN (slo__sro_n714), .A1 (n_11), .A2 (p_1[11]));
NAND3_X1 slo__sro_c477 (.ZN (slo__sro_n713), .A1 (slo__sro_n714), .A2 (slo__sro_n715), .A3 (slo__sro_n716));
XNOR2_X1 slo__sro_c478 (.ZN (slo__sro_n712), .A (p_1[11]), .B (p_0[11]));
XNOR2_X1 slo__sro_c479 (.ZN (p_2[11]), .A (slo__sro_n712), .B (n_11));
NAND2_X1 slo__sro_c491 (.ZN (slo__sro_n736), .A1 (slo__sro_n669), .A2 (p_0[5]));
NAND2_X1 slo__sro_c492 (.ZN (slo__sro_n735), .A1 (p_1[5]), .A2 (slo__sro_n669));
NAND3_X1 slo__sro_c493 (.ZN (slo__sro_n734), .A1 (slo__sro_n735), .A2 (slo__sro_n737), .A3 (slo__sro_n736));
XNOR2_X2 slo__sro_c494 (.ZN (slo__sro_n733), .A (slo__sro_n669), .B (p_0[5]));
XNOR2_X1 slo__sro_c495 (.ZN (p_2[5]), .A (slo__sro_n733), .B (p_1[5]));
XNOR2_X1 slo__mro_c518 (.ZN (p_2[6]), .A (slo__mro_n765), .B (p_1[6]));
XNOR2_X2 CLOCK_slo__mro_c681 (.ZN (p_2[4]), .A (CLOCK_slo__mro_n1112), .B (p_1[4]));
NOR2_X1 CLOCK_slo__sro_c740 (.ZN (CLOCK_slo__sro_n1167), .A1 (p_1[8]), .A2 (p_0[8]));
OAI21_X1 CLOCK_slo__sro_c741 (.ZN (n_9), .A (CLOCK_slo__sro_n1168), .B1 (CLOCK_slo__sro_n1169), .B2 (CLOCK_slo__sro_n1167));
XNOR2_X2 CLOCK_slo__sro_c742 (.ZN (CLOCK_slo__sro_n1166), .A (p_1[8]), .B (p_0[8]));
XNOR2_X1 CLOCK_slo__sro_c743 (.ZN (p_2[8]), .A (CLOCK_slo__sro_n1166), .B (n_8));
INV_X1 CLOCK_slo__sro_c769 (.ZN (CLOCK_slo__sro_n1199), .A (n_24));
NAND2_X1 CLOCK_slo__sro_c770 (.ZN (CLOCK_slo__sro_n1198), .A1 (p_1[24]), .A2 (p_0[24]));
NOR2_X1 CLOCK_slo__sro_c771 (.ZN (CLOCK_slo__sro_n1197), .A1 (p_1[24]), .A2 (p_0[24]));
OAI21_X1 CLOCK_slo__sro_c772 (.ZN (CLOCK_slo__sro_n1196), .A (CLOCK_slo__sro_n1198)
    , .B1 (CLOCK_slo__sro_n1199), .B2 (CLOCK_slo__sro_n1197));
XNOR2_X1 CLOCK_slo__sro_c773 (.ZN (CLOCK_slo__sro_n1195), .A (p_1[24]), .B (p_0[24]));
XNOR2_X1 CLOCK_slo__sro_c774 (.ZN (p_2[24]), .A (n_24), .B (CLOCK_slo__sro_n1195));

endmodule //datapath__0_122

module datapath__0_121 (opt_ipoPP_0, Multiplier, p_0, p_1);

output [31:0] p_1;
input [31:0] Multiplier;
input [31:0] p_0;
input opt_ipoPP_0;
wire slo__sro_n586;
wire CLOCK_slo__sro_n1683;
wire CLOCK_slo__sro_n1291;
wire slo__n1089;
wire n_1;
wire n_2;
wire n_4;
wire n_6;
wire n_7;
wire n_8;
wire n_9;
wire n_10;
wire n_12;
wire n_13;
wire n_16;
wire n_20;
wire n_21;
wire n_22;
wire n_23;
wire n_24;
wire slo__sro_n588;
wire n_27;
wire n_28;
wire n_30;
wire n_32;
wire CLOCK_slo__sro_n1682;
wire n_34;
wire n_33;
wire n_31;
wire slo__sro_n57;
wire slo__sro_n58;
wire slo__sro_n59;
wire slo__sro_n60;
wire CLOCK_slo__n1728;
wire slo__sro_n71;
wire slo__sro_n72;
wire slo__sro_n73;
wire slo__sro_n74;
wire slo__sro_n129;
wire slo__sro_n130;
wire slo__sro_n131;
wire slo__sro_n132;
wire slo__sro_n133;
wire slo__sro_n270;
wire slo__sro_n271;
wire slo__sro_n272;
wire slo__sro_n273;
wire slo__sro_n163;
wire slo__sro_n164;
wire slo__sro_n165;
wire slo__sro_n166;
wire slo__sro_n167;
wire slo__sro_n460;
wire slo__sro_n461;
wire slo__sro_n462;
wire slo__sro_n463;
wire slo__sro_n479;
wire slo__sro_n480;
wire slo__sro_n481;
wire slo__sro_n482;
wire slo__sro_n587;
wire slo__sro_n500;
wire slo__sro_n501;
wire slo__sro_n502;
wire slo__sro_n503;
wire slo__sro_n504;
wire slo__sro_n589;
wire slo__sro_n590;
wire slo__sro_n709;
wire slo__sro_n710;
wire slo__sro_n711;
wire slo__sro_n712;
wire slo__sro_n713;
wire slo__sro_n801;
wire CLOCK_slo__sro_n1292;
wire slo__sro_n803;
wire slo__sro_n987;
wire slo__sro_n988;
wire slo__sro_n989;
wire slo__sro_n990;
wire slo__sro_n991;
wire CLOCK_slo__mro_n1226;
wire CLOCK_slo__sro_n1251;
wire CLOCK_slo__sro_n1293;
wire CLOCK_slo__sro_n1294;
wire CLOCK_slo__sro_n1295;
wire CLOCK_slo__sro_n1308;
wire CLOCK_slo__sro_n1309;
wire CLOCK_slo__sro_n1310;
wire CLOCK_slo__sro_n1311;
wire CLOCK_slo__sro_n1312;
wire CLOCK_slo__sro_n1372;
wire CLOCK_slo__sro_n1373;
wire CLOCK_slo__sro_n1374;
wire CLOCK_slo__sro_n1375;
wire CLOCK_slo__sro_n1398;
wire CLOCK_slo__sro_n1684;
wire CLOCK_slo__sro_n1685;
wire CLOCK_slo__mro_n1692;


INV_X1 i_36 (.ZN (n_34), .A (Multiplier[30]));
INV_X1 i_35 (.ZN (n_33), .A (p_0[30]));
INV_X1 i_34 (.ZN (n_32), .A (n_30));
XNOR2_X1 CLOCK_slo__mro_c1293 (.ZN (CLOCK_slo__mro_n1692), .A (p_0[28]), .B (Multiplier[28]));
XOR2_X1 i_32 (.Z (p_1[31]), .A (Multiplier[31]), .B (n_31));
INV_X1 CLOCK_slo__sro_c1281 (.ZN (CLOCK_slo__sro_n1685), .A (n_30));
XNOR2_X1 i_0 (.ZN (p_1[30]), .A (CLOCK_slo__sro_n1398), .B (n_32));
FA_X1 i_30 (.CO (n_30), .S (p_1[29]), .A (Multiplier[29]), .B (p_0[29]), .CI (slo__sro_n71));
INV_X1 slo__sro_c70 (.ZN (slo__sro_n133), .A (n_2));
NAND2_X1 slo__sro_c454 (.ZN (slo__sro_n589), .A1 (p_0[13]), .A2 (Multiplier[13]));
INV_X1 slo__sro_c369 (.ZN (slo__sro_n482), .A (p_0[27]));
INV_X1 slo__sro_c453 (.ZN (slo__sro_n590), .A (n_13));
OAI21_X1 slo__sro_c456 (.ZN (slo__sro_n587), .A (slo__sro_n589), .B1 (slo__sro_n590), .B2 (slo__sro_n588));
INV_X1 slo__sro_c15 (.ZN (slo__sro_n74), .A (n_28));
FA_X1 i_23 (.CO (n_23), .S (p_1[22]), .A (Multiplier[22]), .B (p_0[22]), .CI (n_22));
FA_X1 i_22 (.CO (n_22), .S (p_1[21]), .A (Multiplier[21]), .B (p_0[21]), .CI (n_21));
FA_X1 i_21 (.CO (n_21), .S (p_1[20]), .A (Multiplier[20]), .B (p_0[20]), .CI (n_20));
FA_X1 i_20 (.CO (n_20), .S (p_1[19]), .A (Multiplier[19]), .B (p_0[19]), .CI (slo__sro_n801));
INV_X2 slo__sro_c744 (.ZN (slo__sro_n991), .A (n_4));
INV_X1 slo__sro_c351 (.ZN (slo__sro_n463), .A (p_0[26]));
INV_X1 CLOCK_slo__sro_c950 (.ZN (CLOCK_slo__sro_n1312), .A (slo__sro_n587));
FA_X1 i_16 (.CO (n_16), .S (p_1[15]), .A (Multiplier[15]), .B (p_0[15]), .CI (CLOCK_slo__sro_n1309));
INV_X1 CLOCK_slo__sro_c1007 (.ZN (CLOCK_slo__sro_n1375), .A (slo__sro_n710));
INV_X1 slo__sro_c548 (.ZN (slo__sro_n713), .A (n_10));
FA_X1 i_13 (.CO (n_13), .S (p_1[12]), .A (Multiplier[12]), .B (p_0[12]), .CI (n_12));
NOR2_X1 CLOCK_slo__sro_c1282 (.ZN (CLOCK_slo__sro_n1684), .A1 (n_33), .A2 (Multiplier[30]));
NAND2_X1 slo__sro_c628 (.ZN (slo__sro_n803), .A1 (p_0[18]), .A2 (Multiplier[18]));
FA_X1 i_10 (.CO (n_10), .S (p_1[9]), .A (Multiplier[9]), .B (p_0[9]), .CI (n_9));
FA_X1 i_9 (.CO (n_9), .S (p_1[8]), .A (Multiplier[8]), .B (p_0[8]), .CI (n_8));
FA_X1 i_8 (.CO (n_8), .S (p_1[7]), .A (Multiplier[7]), .B (p_0[7]), .CI (n_7));
FA_X1 i_7 (.CO (n_7), .S (p_1[6]), .A (Multiplier[6]), .B (p_0[6]), .CI (n_6));
FA_X1 i_6 (.CO (n_6), .S (p_1[5]), .A (Multiplier[5]), .B (p_0[5]), .CI (slo__sro_n988));
OAI21_X1 slo__c822 (.ZN (slo__n1089), .A (slo__sro_n462), .B1 (slo__sro_n463), .B2 (slo__sro_n461));
FA_X1 i_4 (.CO (n_4), .S (p_1[3]), .A (Multiplier[3]), .B (p_0[3]), .CI (slo__sro_n130));
XNOR2_X1 CLOCK_slo__mro_c864 (.ZN (CLOCK_slo__mro_n1226), .A (slo__sro_n164), .B (Multiplier[18]));
FA_X1 i_2 (.CO (n_2), .S (p_1[1]), .A (Multiplier[1]), .B (p_0[1]), .CI (n_1));
HA_X1 i_1 (.CO (n_1), .S (p_1[0]), .A (Multiplier[0]), .B (p_0[0]));
INV_X2 slo__sro_c1 (.ZN (slo__sro_n60), .A (n_23));
NAND2_X1 slo__sro_c2 (.ZN (slo__sro_n59), .A1 (p_0[23]), .A2 (Multiplier[23]));
NOR2_X2 slo__sro_c3 (.ZN (slo__sro_n58), .A1 (p_0[23]), .A2 (Multiplier[23]));
OAI21_X2 slo__sro_c4 (.ZN (n_24), .A (slo__sro_n59), .B1 (slo__sro_n60), .B2 (slo__sro_n58));
XNOR2_X2 slo__sro_c5 (.ZN (slo__sro_n57), .A (p_0[23]), .B (Multiplier[23]));
XNOR2_X2 slo__sro_c6 (.ZN (p_1[23]), .A (slo__sro_n57), .B (n_23));
NAND2_X1 slo__sro_c16 (.ZN (slo__sro_n73), .A1 (p_0[28]), .A2 (Multiplier[28]));
NOR2_X1 slo__sro_c17 (.ZN (slo__sro_n72), .A1 (p_0[28]), .A2 (Multiplier[28]));
OAI21_X1 slo__sro_c18 (.ZN (slo__sro_n71), .A (slo__sro_n73), .B1 (slo__sro_n74), .B2 (slo__sro_n72));
OAI21_X1 CLOCK_slo__c1329 (.ZN (CLOCK_slo__n1728), .A (slo__sro_n481), .B1 (slo__sro_n480), .B2 (slo__sro_n482));
NAND2_X1 slo__sro_c71 (.ZN (slo__sro_n132), .A1 (p_0[2]), .A2 (Multiplier[2]));
NOR2_X1 slo__sro_c72 (.ZN (slo__sro_n131), .A1 (p_0[2]), .A2 (Multiplier[2]));
OAI21_X1 slo__sro_c73 (.ZN (slo__sro_n130), .A (slo__sro_n132), .B1 (slo__sro_n133), .B2 (slo__sro_n131));
XNOR2_X1 slo__sro_c74 (.ZN (slo__sro_n129), .A (p_0[2]), .B (Multiplier[2]));
XNOR2_X1 slo__sro_c75 (.ZN (p_1[2]), .A (slo__sro_n129), .B (n_2));
NAND2_X1 slo__sro_c192 (.ZN (slo__sro_n273), .A1 (slo__sro_n501), .A2 (Multiplier[25]));
NOR2_X2 slo__sro_c193 (.ZN (slo__sro_n272), .A1 (slo__sro_n501), .A2 (Multiplier[25]));
OAI21_X2 slo__sro_c194 (.ZN (slo__sro_n271), .A (slo__sro_n273), .B1 (slo__sro_n272), .B2 (p_0[25]));
XNOR2_X1 slo__sro_c195 (.ZN (slo__sro_n270), .A (slo__sro_n501), .B (Multiplier[25]));
XNOR2_X1 slo__sro_c196 (.ZN (p_1[25]), .A (slo__sro_n270), .B (opt_ipoPP_0));
INV_X1 slo__sro_c99 (.ZN (slo__sro_n167), .A (CLOCK_slo__sro_n1292));
NAND2_X1 slo__sro_c100 (.ZN (slo__sro_n166), .A1 (p_0[17]), .A2 (Multiplier[17]));
NOR2_X1 slo__sro_c101 (.ZN (slo__sro_n165), .A1 (p_0[17]), .A2 (Multiplier[17]));
OAI21_X1 slo__sro_c102 (.ZN (slo__sro_n164), .A (slo__sro_n166), .B1 (slo__sro_n167), .B2 (slo__sro_n165));
XNOR2_X1 slo__sro_c103 (.ZN (slo__sro_n163), .A (p_0[17]), .B (Multiplier[17]));
XNOR2_X1 slo__sro_c104 (.ZN (p_1[17]), .A (CLOCK_slo__sro_n1292), .B (slo__sro_n163));
NAND2_X1 slo__sro_c352 (.ZN (slo__sro_n462), .A1 (slo__sro_n271), .A2 (Multiplier[26]));
NOR2_X1 CLOCK_slo__sro_c938 (.ZN (CLOCK_slo__sro_n1293), .A1 (p_0[16]), .A2 (Multiplier[16]));
OAI21_X2 slo__sro_c354 (.ZN (n_27), .A (slo__sro_n462), .B1 (slo__sro_n463), .B2 (slo__sro_n461));
XNOR2_X2 slo__sro_c355 (.ZN (slo__sro_n460), .A (slo__sro_n271), .B (Multiplier[26]));
XNOR2_X2 slo__sro_c356 (.ZN (p_1[26]), .A (slo__sro_n460), .B (p_0[26]));
NAND2_X1 slo__sro_c370 (.ZN (slo__sro_n481), .A1 (n_27), .A2 (Multiplier[27]));
NOR2_X1 slo__sro_c371 (.ZN (slo__sro_n480), .A1 (n_27), .A2 (Multiplier[27]));
OAI21_X1 slo__sro_c372 (.ZN (n_28), .A (slo__sro_n481), .B1 (slo__sro_n480), .B2 (slo__sro_n482));
XNOR2_X1 slo__sro_c373 (.ZN (slo__sro_n479), .A (slo__n1089), .B (Multiplier[27]));
XNOR2_X1 slo__sro_c374 (.ZN (p_1[27]), .A (slo__sro_n479), .B (p_0[27]));
NOR2_X1 slo__sro_c455 (.ZN (slo__sro_n588), .A1 (p_0[13]), .A2 (Multiplier[13]));
INV_X2 slo__sro_c389 (.ZN (slo__sro_n504), .A (n_24));
NAND2_X1 slo__sro_c390 (.ZN (slo__sro_n503), .A1 (p_0[24]), .A2 (Multiplier[24]));
NOR2_X1 slo__sro_c391 (.ZN (slo__sro_n502), .A1 (p_0[24]), .A2 (Multiplier[24]));
OAI21_X2 slo__sro_c392 (.ZN (slo__sro_n501), .A (slo__sro_n503), .B1 (slo__sro_n504), .B2 (slo__sro_n502));
XNOR2_X1 slo__sro_c393 (.ZN (slo__sro_n500), .A (p_0[24]), .B (Multiplier[24]));
XNOR2_X1 slo__sro_c394 (.ZN (p_1[24]), .A (n_24), .B (slo__sro_n500));
XNOR2_X1 slo__sro_c457 (.ZN (slo__sro_n586), .A (p_0[13]), .B (Multiplier[13]));
XNOR2_X1 slo__sro_c458 (.ZN (p_1[13]), .A (n_13), .B (slo__sro_n586));
NAND2_X1 slo__sro_c549 (.ZN (slo__sro_n712), .A1 (p_0[10]), .A2 (Multiplier[10]));
NOR2_X1 slo__sro_c550 (.ZN (slo__sro_n711), .A1 (p_0[10]), .A2 (Multiplier[10]));
OAI21_X1 slo__sro_c551 (.ZN (slo__sro_n710), .A (slo__sro_n712), .B1 (slo__sro_n711), .B2 (slo__sro_n713));
XNOR2_X1 slo__sro_c552 (.ZN (slo__sro_n709), .A (p_0[10]), .B (Multiplier[10]));
XNOR2_X1 slo__sro_c553 (.ZN (p_1[10]), .A (slo__sro_n709), .B (n_10));
OAI21_X1 CLOCK_slo__sro_c939 (.ZN (CLOCK_slo__sro_n1292), .A (CLOCK_slo__sro_n1294)
    , .B1 (CLOCK_slo__sro_n1295), .B2 (CLOCK_slo__sro_n1293));
NAND2_X1 slo__sro_c630 (.ZN (slo__sro_n801), .A1 (CLOCK_slo__sro_n1251), .A2 (slo__sro_n803));
INV_X1 CLOCK_slo__sro_c936 (.ZN (CLOCK_slo__sro_n1295), .A (n_16));
NAND2_X1 CLOCK_slo__sro_c937 (.ZN (CLOCK_slo__sro_n1294), .A1 (p_0[16]), .A2 (Multiplier[16]));
NAND2_X1 slo__sro_c745 (.ZN (slo__sro_n990), .A1 (p_0[4]), .A2 (Multiplier[4]));
NOR2_X1 slo__sro_c746 (.ZN (slo__sro_n989), .A1 (p_0[4]), .A2 (Multiplier[4]));
OAI21_X2 slo__sro_c747 (.ZN (slo__sro_n988), .A (slo__sro_n990), .B1 (slo__sro_n991), .B2 (slo__sro_n989));
XNOR2_X1 slo__sro_c748 (.ZN (slo__sro_n987), .A (p_0[4]), .B (Multiplier[4]));
XNOR2_X1 slo__sro_c749 (.ZN (p_1[4]), .A (slo__sro_n987), .B (n_4));
XNOR2_X1 CLOCK_slo__mro_c865 (.ZN (p_1[18]), .A (CLOCK_slo__mro_n1226), .B (p_0[18]));
NOR2_X2 CLOCK_slo__mro_c877 (.ZN (slo__sro_n461), .A1 (slo__sro_n271), .A2 (Multiplier[26]));
OAI21_X1 CLOCK_slo__sro_c902 (.ZN (CLOCK_slo__sro_n1251), .A (slo__sro_n164), .B1 (p_0[18]), .B2 (Multiplier[18]));
XNOR2_X1 CLOCK_slo__sro_c940 (.ZN (CLOCK_slo__sro_n1291), .A (p_0[16]), .B (Multiplier[16]));
XNOR2_X1 CLOCK_slo__sro_c941 (.ZN (p_1[16]), .A (CLOCK_slo__sro_n1291), .B (n_16));
NAND2_X1 CLOCK_slo__sro_c951 (.ZN (CLOCK_slo__sro_n1311), .A1 (p_0[14]), .A2 (Multiplier[14]));
NOR2_X1 CLOCK_slo__sro_c952 (.ZN (CLOCK_slo__sro_n1310), .A1 (p_0[14]), .A2 (Multiplier[14]));
OAI21_X1 CLOCK_slo__sro_c953 (.ZN (CLOCK_slo__sro_n1309), .A (CLOCK_slo__sro_n1311)
    , .B1 (CLOCK_slo__sro_n1312), .B2 (CLOCK_slo__sro_n1310));
XNOR2_X2 CLOCK_slo__sro_c954 (.ZN (CLOCK_slo__sro_n1308), .A (p_0[14]), .B (Multiplier[14]));
XNOR2_X1 CLOCK_slo__sro_c955 (.ZN (p_1[14]), .A (slo__sro_n587), .B (CLOCK_slo__sro_n1308));
NAND2_X1 CLOCK_slo__sro_c1008 (.ZN (CLOCK_slo__sro_n1374), .A1 (p_0[11]), .A2 (Multiplier[11]));
NOR2_X1 CLOCK_slo__sro_c1009 (.ZN (CLOCK_slo__sro_n1373), .A1 (p_0[11]), .A2 (Multiplier[11]));
OAI21_X1 CLOCK_slo__sro_c1010 (.ZN (n_12), .A (CLOCK_slo__sro_n1374), .B1 (CLOCK_slo__sro_n1375), .B2 (CLOCK_slo__sro_n1373));
XNOR2_X1 CLOCK_slo__sro_c1011 (.ZN (CLOCK_slo__sro_n1372), .A (p_0[11]), .B (Multiplier[11]));
XNOR2_X1 CLOCK_slo__sro_c1012 (.ZN (p_1[11]), .A (CLOCK_slo__sro_n1372), .B (slo__sro_n710));
OAI22_X1 CLOCK_slo__sro_c1040 (.ZN (CLOCK_slo__sro_n1398), .A1 (n_33), .A2 (Multiplier[30])
    , .B1 (p_0[30]), .B2 (n_34));
NAND2_X1 CLOCK_slo__sro_c1283 (.ZN (CLOCK_slo__sro_n1683), .A1 (CLOCK_slo__sro_n1684), .A2 (CLOCK_slo__sro_n1685));
OR2_X1 CLOCK_slo__sro_c1284 (.ZN (CLOCK_slo__sro_n1682), .A1 (p_0[30]), .A2 (n_34));
OAI21_X1 CLOCK_slo__sro_c1285 (.ZN (n_31), .A (CLOCK_slo__sro_n1683), .B1 (n_32), .B2 (CLOCK_slo__sro_n1682));
XNOR2_X1 CLOCK_slo__mro_c1294 (.ZN (p_1[28]), .A (CLOCK_slo__mro_n1692), .B (CLOCK_slo__n1728));

endmodule //datapath__0_121

module datapath__0_117 (p_0, p_1, p_2);

output [31:0] p_2;
input [31:0] p_0;
input [31:0] p_1;
wire CLOCK_slo__sro_n1207;
wire n_1;
wire n_2;
wire n_3;
wire n_4;
wire n_5;
wire n_6;
wire n_7;
wire n_8;
wire n_9;
wire n_10;
wire n_11;
wire n_12;
wire n_13;
wire n_14;
wire n_17;
wire n_18;
wire n_19;
wire n_20;
wire n_21;
wire n_22;
wire n_23;
wire n_24;
wire n_25;
wire n_27;
wire n_28;
wire n_32;
wire n_0;
wire n_34;
wire n_33;
wire n_31;
wire slo__sro_n65;
wire slo__sro_n66;
wire slo__sro_n67;
wire slo__sro_n68;
wire slo__sro_n147;
wire slo__sro_n148;
wire slo__sro_n149;
wire slo__sro_n150;
wire slo__sro_n253;
wire slo__sro_n254;
wire slo__sro_n255;
wire slo__sro_n256;
wire slo__sro_n176;
wire slo__sro_n177;
wire slo__sro_n178;
wire slo__sro_n179;
wire slo__sro_n180;
wire slo__sro_n338;
wire slo__sro_n339;
wire slo__sro_n340;
wire slo__sro_n341;
wire slo__sro_n342;
wire slo__sro_n618;
wire slo__sro_n619;
wire slo__sro_n620;
wire slo__sro_n621;
wire slo__sro_n622;
wire CLOCK_slo__sro_n964;
wire CLOCK_slo__sro_n965;
wire CLOCK_slo__sro_n966;
wire CLOCK_slo__sro_n967;
wire CLOCK_slo__sro_n979;
wire CLOCK_slo__sro_n980;
wire CLOCK_slo__sro_n981;
wire CLOCK_slo__sro_n982;
wire CLOCK_slo__sro_n993;
wire slo__sro_n323;
wire slo__sro_n324;
wire slo__sro_n325;
wire slo__sro_n326;
wire CLOCK_slo__sro_n994;
wire CLOCK_slo__sro_n995;
wire CLOCK_slo__sro_n996;
wire CLOCK_slo__sro_n997;
wire CLOCK_slo__sro_n1039;
wire CLOCK_slo__sro_n1040;
wire CLOCK_slo__sro_n1041;
wire CLOCK_slo__sro_n1042;
wire CLOCK_slo__sro_n1056;
wire CLOCK_slo__sro_n1057;
wire CLOCK_slo__sro_n1058;
wire CLOCK_slo__sro_n1059;
wire CLOCK_slo__sro_n1204;
wire CLOCK_slo__sro_n1205;
wire CLOCK_slo__sro_n1206;
wire CLOCK_slo__sro_n1097;
wire CLOCK_slo__sro_n1098;
wire CLOCK_slo__sro_n1099;
wire CLOCK_slo__sro_n1100;
wire CLOCK_slo__sro_n1208;


INV_X1 i_36 (.ZN (n_34), .A (p_0[30]));
INV_X1 i_35 (.ZN (n_33), .A (p_1[30]));
INV_X1 i_34 (.ZN (n_32), .A (slo__sro_n177));
NAND2_X1 CLOCK_slo__sro_c667 (.ZN (CLOCK_slo__sro_n996), .A1 (p_1[14]), .A2 (p_0[14]));
XOR2_X1 i_32 (.Z (p_2[31]), .A (p_0[31]), .B (n_31));
OAI22_X1 i_31 (.ZN (n_0), .A1 (n_34), .A2 (p_1[30]), .B1 (n_33), .B2 (p_0[30]));
XNOR2_X1 i_0 (.ZN (p_2[30]), .A (n_32), .B (n_0));
NAND2_X1 slo__sro_c238 (.ZN (slo__sro_n341), .A1 (p_1[28]), .A2 (p_0[28]));
XNOR2_X1 CLOCK_slo__sro_c859 (.ZN (p_2[25]), .A (CLOCK_slo__sro_n1204), .B (n_25));
FA_X1 i_27 (.CO (n_27), .S (p_2[26]), .A (p_0[26]), .B (p_1[26]), .CI (CLOCK_slo__sro_n1205));
FA_X1 i_25 (.CO (n_25), .S (p_2[24]), .A (p_0[24]), .B (p_1[24]), .CI (n_24));
FA_X1 i_24 (.CO (n_24), .S (p_2[23]), .A (p_0[23]), .B (p_1[23]), .CI (n_23));
INV_X1 slo__sro_c237 (.ZN (slo__sro_n342), .A (n_28));
FA_X1 i_22 (.CO (n_22), .S (p_2[21]), .A (p_0[21]), .B (p_1[21]), .CI (n_21));
FA_X1 i_21 (.CO (n_21), .S (p_2[20]), .A (p_0[20]), .B (p_1[20]), .CI (n_20));
FA_X1 i_20 (.CO (n_20), .S (p_2[19]), .A (p_0[19]), .B (p_1[19]), .CI (n_19));
INV_X1 slo__sro_c82 (.ZN (slo__sro_n150), .A (n_3));
FA_X1 i_18 (.CO (n_18), .S (p_2[17]), .A (p_0[17]), .B (p_1[17]), .CI (n_17));
FA_X1 i_17 (.CO (n_17), .S (p_2[16]), .A (p_0[16]), .B (p_1[16]), .CI (slo__sro_n619));
INV_X1 CLOCK_slo__sro_c628 (.ZN (CLOCK_slo__sro_n967), .A (n_5));
INV_X1 CLOCK_slo__sro_c708 (.ZN (CLOCK_slo__sro_n1042), .A (n_11));
FA_X1 i_14 (.CO (n_14), .S (p_2[13]), .A (p_0[13]), .B (p_1[13]), .CI (n_13));
FA_X1 i_13 (.CO (n_13), .S (p_2[12]), .A (p_0[12]), .B (p_1[12]), .CI (n_12));
INV_X2 CLOCK_slo__sro_c724 (.ZN (CLOCK_slo__sro_n1059), .A (n_10));
OAI21_X2 CLOCK_slo__sro_c837 (.ZN (n_4), .A (slo__sro_n149), .B1 (slo__sro_n148), .B2 (slo__sro_n150));
FA_X1 i_10 (.CO (n_10), .S (p_2[9]), .A (p_0[9]), .B (p_1[9]), .CI (n_9));
FA_X1 i_9 (.CO (n_9), .S (p_2[8]), .A (p_0[8]), .B (p_1[8]), .CI (n_8));
FA_X1 i_8 (.CO (n_8), .S (p_2[7]), .A (p_0[7]), .B (p_1[7]), .CI (n_7));
FA_X1 i_7 (.CO (n_7), .S (p_2[6]), .A (p_0[6]), .B (p_1[6]), .CI (n_6));
INV_X1 CLOCK_slo__sro_c666 (.ZN (CLOCK_slo__sro_n997), .A (n_14));
FA_X1 i_5 (.CO (n_5), .S (p_2[4]), .A (p_0[4]), .B (p_1[4]), .CI (n_4));
INV_X1 slo__sro_c155 (.ZN (slo__sro_n256), .A (n_22));
FA_X1 i_3 (.CO (n_3), .S (p_2[2]), .A (p_0[2]), .B (p_1[2]), .CI (n_2));
OAI21_X2 CLOCK_slo__sro_c669 (.ZN (CLOCK_slo__sro_n994), .A (CLOCK_slo__sro_n996)
    , .B1 (CLOCK_slo__sro_n997), .B2 (CLOCK_slo__sro_n995));
HA_X1 i_1 (.CO (n_1), .S (p_2[0]), .A (p_0[0]), .B (p_1[0]));
INV_X1 slo__sro_c3 (.ZN (slo__sro_n68), .A (n_18));
NAND2_X1 slo__sro_c4 (.ZN (slo__sro_n67), .A1 (p_1[18]), .A2 (p_0[18]));
NOR2_X1 slo__sro_c5 (.ZN (slo__sro_n66), .A1 (p_1[18]), .A2 (p_0[18]));
OAI21_X1 slo__sro_c6 (.ZN (n_19), .A (slo__sro_n67), .B1 (slo__sro_n68), .B2 (slo__sro_n66));
XNOR2_X1 slo__sro_c7 (.ZN (slo__sro_n65), .A (p_1[18]), .B (p_0[18]));
XNOR2_X1 slo__sro_c8 (.ZN (p_2[18]), .A (slo__sro_n65), .B (n_18));
NAND2_X1 slo__sro_c83 (.ZN (slo__sro_n149), .A1 (p_1[3]), .A2 (p_0[3]));
NOR2_X1 slo__sro_c84 (.ZN (slo__sro_n148), .A1 (p_1[3]), .A2 (p_0[3]));
XNOR2_X1 slo__sro_c86 (.ZN (slo__sro_n147), .A (p_1[3]), .B (p_0[3]));
XNOR2_X1 slo__sro_c87 (.ZN (p_2[3]), .A (slo__sro_n147), .B (n_3));
NAND2_X1 slo__sro_c156 (.ZN (slo__sro_n255), .A1 (p_1[22]), .A2 (p_0[22]));
NOR2_X1 slo__sro_c157 (.ZN (slo__sro_n254), .A1 (p_1[22]), .A2 (p_0[22]));
OAI21_X1 slo__sro_c158 (.ZN (n_23), .A (slo__sro_n255), .B1 (slo__sro_n256), .B2 (slo__sro_n254));
XNOR2_X1 slo__sro_c159 (.ZN (slo__sro_n253), .A (p_1[22]), .B (p_0[22]));
XNOR2_X1 slo__sro_c160 (.ZN (p_2[22]), .A (n_22), .B (slo__sro_n253));
INV_X1 slo__sro_c113 (.ZN (slo__sro_n180), .A (slo__sro_n339));
NAND2_X1 slo__sro_c114 (.ZN (slo__sro_n179), .A1 (p_1[29]), .A2 (p_0[29]));
NOR2_X1 slo__sro_c115 (.ZN (slo__sro_n178), .A1 (p_1[29]), .A2 (p_0[29]));
OAI21_X1 slo__sro_c116 (.ZN (slo__sro_n177), .A (slo__sro_n179), .B1 (slo__sro_n180), .B2 (slo__sro_n178));
XNOR2_X1 slo__sro_c117 (.ZN (slo__sro_n176), .A (p_1[29]), .B (p_0[29]));
XNOR2_X1 slo__sro_c118 (.ZN (p_2[29]), .A (slo__sro_n339), .B (slo__sro_n176));
NOR2_X1 slo__sro_c239 (.ZN (slo__sro_n340), .A1 (p_1[28]), .A2 (p_0[28]));
OAI21_X1 slo__sro_c240 (.ZN (slo__sro_n339), .A (slo__sro_n341), .B1 (slo__sro_n342), .B2 (slo__sro_n340));
XNOR2_X1 slo__sro_c241 (.ZN (slo__sro_n338), .A (p_1[28]), .B (p_0[28]));
XNOR2_X1 slo__sro_c242 (.ZN (p_2[28]), .A (slo__sro_n338), .B (n_28));
INV_X1 slo__sro_c441 (.ZN (slo__sro_n622), .A (CLOCK_slo__sro_n994));
NAND2_X1 slo__sro_c442 (.ZN (slo__sro_n621), .A1 (p_1[15]), .A2 (p_0[15]));
NOR2_X1 slo__sro_c443 (.ZN (slo__sro_n620), .A1 (p_1[15]), .A2 (p_0[15]));
OAI21_X1 slo__sro_c444 (.ZN (slo__sro_n619), .A (slo__sro_n621), .B1 (slo__sro_n622), .B2 (slo__sro_n620));
XNOR2_X1 slo__sro_c445 (.ZN (slo__sro_n618), .A (p_1[15]), .B (p_0[15]));
XNOR2_X1 slo__sro_c446 (.ZN (p_2[15]), .A (slo__sro_n618), .B (CLOCK_slo__sro_n994));
NAND2_X1 CLOCK_slo__sro_c629 (.ZN (CLOCK_slo__sro_n966), .A1 (p_1[5]), .A2 (p_0[5]));
NOR2_X1 CLOCK_slo__sro_c630 (.ZN (CLOCK_slo__sro_n965), .A1 (p_1[5]), .A2 (p_0[5]));
OAI21_X2 CLOCK_slo__sro_c631 (.ZN (n_6), .A (CLOCK_slo__sro_n966), .B1 (CLOCK_slo__sro_n967), .B2 (CLOCK_slo__sro_n965));
XNOR2_X2 CLOCK_slo__sro_c632 (.ZN (CLOCK_slo__sro_n964), .A (p_1[5]), .B (p_0[5]));
XNOR2_X2 CLOCK_slo__sro_c633 (.ZN (p_2[5]), .A (CLOCK_slo__sro_n964), .B (n_5));
INV_X1 CLOCK_slo__sro_c649 (.ZN (CLOCK_slo__sro_n982), .A (n_34));
INV_X1 CLOCK_slo__sro_c650 (.ZN (CLOCK_slo__sro_n981), .A (p_1[30]));
OR2_X1 CLOCK_slo__sro_c651 (.ZN (CLOCK_slo__sro_n980), .A1 (n_33), .A2 (p_0[30]));
NAND2_X1 CLOCK_slo__sro_c652 (.ZN (CLOCK_slo__sro_n979), .A1 (CLOCK_slo__sro_n981), .A2 (CLOCK_slo__sro_n982));
OAI22_X1 CLOCK_slo__sro_c653 (.ZN (n_31), .A1 (n_32), .A2 (CLOCK_slo__sro_n979), .B1 (CLOCK_slo__sro_n980), .B2 (slo__sro_n177));
NOR2_X1 CLOCK_slo__sro_c668 (.ZN (CLOCK_slo__sro_n995), .A1 (p_1[14]), .A2 (p_0[14]));
INV_X2 slo__sro_c221 (.ZN (slo__sro_n326), .A (p_1[1]));
NAND2_X1 slo__sro_c222 (.ZN (slo__sro_n325), .A1 (n_1), .A2 (p_0[1]));
NOR2_X1 slo__sro_c223 (.ZN (slo__sro_n324), .A1 (n_1), .A2 (p_0[1]));
OAI21_X2 slo__sro_c224 (.ZN (n_2), .A (slo__sro_n325), .B1 (slo__sro_n326), .B2 (slo__sro_n324));
XNOR2_X1 slo__sro_c225 (.ZN (slo__sro_n323), .A (n_1), .B (p_0[1]));
XNOR2_X1 slo__sro_c226 (.ZN (p_2[1]), .A (slo__sro_n323), .B (p_1[1]));
XNOR2_X1 CLOCK_slo__sro_c670 (.ZN (CLOCK_slo__sro_n993), .A (p_1[14]), .B (p_0[14]));
XNOR2_X1 CLOCK_slo__sro_c671 (.ZN (p_2[14]), .A (n_14), .B (CLOCK_slo__sro_n993));
NAND2_X1 CLOCK_slo__sro_c709 (.ZN (CLOCK_slo__sro_n1041), .A1 (p_1[11]), .A2 (p_0[11]));
NOR2_X1 CLOCK_slo__sro_c710 (.ZN (CLOCK_slo__sro_n1040), .A1 (p_1[11]), .A2 (p_0[11]));
OAI21_X1 CLOCK_slo__sro_c711 (.ZN (n_12), .A (CLOCK_slo__sro_n1041), .B1 (CLOCK_slo__sro_n1042), .B2 (CLOCK_slo__sro_n1040));
XNOR2_X1 CLOCK_slo__sro_c712 (.ZN (CLOCK_slo__sro_n1039), .A (p_1[11]), .B (p_0[11]));
XNOR2_X1 CLOCK_slo__sro_c713 (.ZN (p_2[11]), .A (n_11), .B (CLOCK_slo__sro_n1039));
NAND2_X1 CLOCK_slo__sro_c725 (.ZN (CLOCK_slo__sro_n1058), .A1 (p_1[10]), .A2 (p_0[10]));
NOR2_X1 CLOCK_slo__sro_c726 (.ZN (CLOCK_slo__sro_n1057), .A1 (p_1[10]), .A2 (p_0[10]));
OAI21_X2 CLOCK_slo__sro_c727 (.ZN (n_11), .A (CLOCK_slo__sro_n1058), .B1 (CLOCK_slo__sro_n1059), .B2 (CLOCK_slo__sro_n1057));
XNOR2_X1 CLOCK_slo__sro_c728 (.ZN (CLOCK_slo__sro_n1056), .A (p_1[10]), .B (p_0[10]));
XNOR2_X1 CLOCK_slo__sro_c729 (.ZN (p_2[10]), .A (CLOCK_slo__sro_n1056), .B (n_10));
INV_X1 CLOCK_slo__sro_c854 (.ZN (CLOCK_slo__sro_n1208), .A (n_25));
NAND2_X1 CLOCK_slo__sro_c855 (.ZN (CLOCK_slo__sro_n1207), .A1 (p_1[25]), .A2 (p_0[25]));
NOR2_X1 CLOCK_slo__sro_c856 (.ZN (CLOCK_slo__sro_n1206), .A1 (p_1[25]), .A2 (p_0[25]));
OAI21_X1 CLOCK_slo__sro_c857 (.ZN (CLOCK_slo__sro_n1205), .A (CLOCK_slo__sro_n1207)
    , .B1 (CLOCK_slo__sro_n1206), .B2 (CLOCK_slo__sro_n1208));
XNOR2_X1 CLOCK_slo__sro_c858 (.ZN (CLOCK_slo__sro_n1204), .A (p_1[25]), .B (p_0[25]));
INV_X1 CLOCK_slo__sro_c775 (.ZN (CLOCK_slo__sro_n1100), .A (n_27));
NAND2_X1 CLOCK_slo__sro_c776 (.ZN (CLOCK_slo__sro_n1099), .A1 (p_1[27]), .A2 (p_0[27]));
NOR2_X1 CLOCK_slo__sro_c777 (.ZN (CLOCK_slo__sro_n1098), .A1 (p_1[27]), .A2 (p_0[27]));
OAI21_X1 CLOCK_slo__sro_c778 (.ZN (n_28), .A (CLOCK_slo__sro_n1099), .B1 (CLOCK_slo__sro_n1100), .B2 (CLOCK_slo__sro_n1098));
XNOR2_X1 CLOCK_slo__sro_c779 (.ZN (CLOCK_slo__sro_n1097), .A (p_1[27]), .B (p_0[27]));
XNOR2_X1 CLOCK_slo__sro_c780 (.ZN (p_2[27]), .A (CLOCK_slo__sro_n1097), .B (n_27));

endmodule //datapath__0_117

module datapath__0_116 (opt_ipoPP_2, Multiplier, p_0, p_1);

output [31:0] p_1;
input [31:0] Multiplier;
input [31:0] p_0;
input opt_ipoPP_2;
wire slo__sro_n556;
wire CLOCK_slo__sro_n1457;
wire n_1;
wire n_2;
wire n_3;
wire n_4;
wire n_5;
wire n_6;
wire n_7;
wire n_8;
wire n_9;
wire n_12;
wire n_14;
wire n_15;
wire n_17;
wire n_18;
wire n_19;
wire n_22;
wire n_23;
wire n_24;
wire n_25;
wire n_26;
wire n_27;
wire slo__sro_n557;
wire n_30;
wire n_32;
wire n_0;
wire n_34;
wire slo__sro_n743;
wire n_31;
wire slo__sro_n129;
wire slo__sro_n130;
wire slo__sro_n131;
wire slo__sro_n132;
wire slo__sro_n133;
wire slo__sro_n176;
wire slo__sro_n177;
wire slo__sro_n178;
wire slo__sro_n179;
wire slo__sro_n180;
wire slo__sro_n207;
wire slo__sro_n208;
wire slo__sro_n209;
wire slo__sro_n210;
wire slo__sro_n332;
wire slo__sro_n333;
wire slo__sro_n334;
wire slo__sro_n335;
wire slo__sro_n336;
wire CLOCK_slo__mro_n1800;
wire slo__sro_n352;
wire slo__sro_n353;
wire slo__sro_n354;
wire slo__sro_n454;
wire slo__sro_n455;
wire slo__sro_n456;
wire slo__sro_n457;
wire slo__sro_n458;
wire slo__sro_n558;
wire slo__sro_n559;
wire slo__sro_n560;
wire slo__sro_n618;
wire slo__sro_n619;
wire slo__sro_n620;
wire slo__sro_n621;
wire slo__sro_n637;
wire slo__sro_n638;
wire slo__sro_n639;
wire slo__sro_n742;
wire slo__sro_n744;
wire slo__sro_n745;
wire slo__sro_n746;
wire CLOCK_slo__sro_n1456;
wire CLOCK_slo__sro_n1458;
wire CLOCK_slo__sro_n1459;
wire CLOCK_slo__sro_n1460;
wire CLOCK_slo__sro_n1475;
wire CLOCK_slo__sro_n1476;
wire CLOCK_slo__sro_n1477;
wire CLOCK_slo__sro_n1478;
wire CLOCK_slo__sro_n1492;
wire CLOCK_slo__sro_n1493;
wire slo__sro_n543;
wire slo__sro_n544;
wire slo__sro_n545;
wire slo__sro_n546;
wire CLOCK_slo__sro_n1494;
wire CLOCK_slo__sro_n1495;
wire CLOCK_slo__sro_n1496;


INV_X1 i_36 (.ZN (n_34), .A (Multiplier[30]));
INV_X1 slo__sro_c577 (.ZN (slo__sro_n746), .A (n_12));
INV_X1 i_34 (.ZN (n_32), .A (n_30));
OAI33_X1 i_33 (.ZN (n_31), .A1 (n_32), .A2 (opt_ipoPP_2), .A3 (n_34), .B1 (n_30), .B2 (p_0[30]), .B3 (Multiplier[30]));
XOR2_X1 i_32 (.Z (p_1[31]), .A (Multiplier[31]), .B (n_31));
OAI22_X1 i_31 (.ZN (n_0), .A1 (opt_ipoPP_2), .A2 (n_34), .B1 (Multiplier[30]), .B2 (p_0[30]));
XNOR2_X1 i_0 (.ZN (p_1[30]), .A (n_32), .B (n_0));
INV_X1 slo__sro_c421 (.ZN (slo__sro_n560), .A (n_15));
NOR2_X1 slo__sro_c423 (.ZN (slo__sro_n558), .A1 (p_0[15]), .A2 (Multiplier[15]));
INV_X1 slo__sro_c255 (.ZN (slo__sro_n354), .A (n_25));
NAND2_X1 slo__sro_c578 (.ZN (slo__sro_n745), .A1 (p_0[12]), .A2 (Multiplier[12]));
NAND2_X1 slo__sro_c422 (.ZN (slo__sro_n559), .A1 (p_0[15]), .A2 (Multiplier[15]));
FA_X1 i_25 (.CO (n_25), .S (p_1[24]), .A (Multiplier[24]), .B (p_0[24]), .CI (n_24));
FA_X1 i_24 (.CO (n_24), .S (p_1[23]), .A (Multiplier[23]), .B (p_0[23]), .CI (n_23));
FA_X1 i_23 (.CO (n_23), .S (p_1[22]), .A (Multiplier[22]), .B (p_0[22]), .CI (n_22));
FA_X1 i_22 (.CO (n_22), .S (p_1[21]), .A (Multiplier[21]), .B (p_0[21]), .CI (slo__sro_n130));
INV_X1 slo__sro_c106 (.ZN (slo__sro_n180), .A (n_9));
FA_X1 i_19 (.CO (n_19), .S (p_1[18]), .A (Multiplier[18]), .B (p_0[18]), .CI (n_18));
FA_X1 i_18 (.CO (n_18), .S (p_1[17]), .A (Multiplier[17]), .B (p_0[17]), .CI (n_17));
FA_X1 i_17 (.CO (n_17), .S (p_1[16]), .A (Multiplier[16]), .B (p_0[16]), .CI (slo__sro_n557));
INV_X1 slo__sro_c476 (.ZN (slo__sro_n621), .A (n_14));
NAND2_X1 slo__sro_c497 (.ZN (slo__sro_n639), .A1 (n_26), .A2 (Multiplier[26]));
FA_X1 i_14 (.CO (n_14), .S (p_1[13]), .A (Multiplier[13]), .B (p_0[13]), .CI (slo__sro_n743));
NOR2_X1 CLOCK_slo__sro_c1127 (.ZN (CLOCK_slo__sro_n1458), .A1 (p_0[10]), .A2 (Multiplier[10]));
FA_X1 i_12 (.CO (n_12), .S (p_1[11]), .A (Multiplier[11]), .B (p_0[11]), .CI (CLOCK_slo__sro_n1457));
INV_X2 CLOCK_slo__sro_c1142 (.ZN (CLOCK_slo__sro_n1478), .A (n_7));
INV_X1 slo__sro_c135 (.ZN (slo__sro_n210), .A (slo__sro_n455));
FA_X1 i_9 (.CO (n_9), .S (p_1[8]), .A (Multiplier[8]), .B (p_0[8]), .CI (n_8));
INV_X1 CLOCK_slo__sro_c1158 (.ZN (CLOCK_slo__sro_n1496), .A (n_19));
FA_X1 i_7 (.CO (n_7), .S (p_1[6]), .A (Multiplier[6]), .B (p_0[6]), .CI (n_6));
FA_X1 i_6 (.CO (n_6), .S (p_1[5]), .A (Multiplier[5]), .B (p_0[5]), .CI (n_5));
FA_X1 i_5 (.CO (n_5), .S (p_1[4]), .A (Multiplier[4]), .B (p_0[4]), .CI (n_4));
FA_X1 i_4 (.CO (n_4), .S (p_1[3]), .A (Multiplier[3]), .B (p_0[3]), .CI (n_3));
FA_X1 i_3 (.CO (n_3), .S (p_1[2]), .A (Multiplier[2]), .B (p_0[2]), .CI (n_2));
NOR2_X1 CLOCK_slo__sro_c1160 (.ZN (CLOCK_slo__sro_n1494), .A1 (p_0[19]), .A2 (Multiplier[19]));
HA_X1 i_1 (.CO (n_1), .S (p_1[0]), .A (Multiplier[0]), .B (p_0[0]));
INV_X2 slo__sro_c66 (.ZN (slo__sro_n133), .A (CLOCK_slo__sro_n1493));
NAND2_X1 slo__sro_c67 (.ZN (slo__sro_n132), .A1 (p_0[20]), .A2 (Multiplier[20]));
NOR2_X2 slo__sro_c68 (.ZN (slo__sro_n131), .A1 (p_0[20]), .A2 (Multiplier[20]));
OAI21_X1 slo__sro_c69 (.ZN (slo__sro_n130), .A (slo__sro_n132), .B1 (slo__sro_n133), .B2 (slo__sro_n131));
XNOR2_X1 slo__sro_c70 (.ZN (slo__sro_n129), .A (p_0[20]), .B (Multiplier[20]));
XNOR2_X1 slo__sro_c71 (.ZN (p_1[20]), .A (CLOCK_slo__sro_n1493), .B (slo__sro_n129));
NAND2_X1 slo__sro_c107 (.ZN (slo__sro_n179), .A1 (p_0[9]), .A2 (Multiplier[9]));
NOR2_X1 slo__sro_c108 (.ZN (slo__sro_n178), .A1 (p_0[9]), .A2 (Multiplier[9]));
OAI21_X1 slo__sro_c109 (.ZN (slo__sro_n177), .A (slo__sro_n179), .B1 (slo__sro_n180), .B2 (slo__sro_n178));
XNOR2_X1 slo__sro_c110 (.ZN (slo__sro_n176), .A (p_0[9]), .B (Multiplier[9]));
XNOR2_X1 slo__sro_c111 (.ZN (p_1[9]), .A (n_9), .B (slo__sro_n176));
NAND2_X1 slo__sro_c136 (.ZN (slo__sro_n209), .A1 (p_0[29]), .A2 (Multiplier[29]));
NOR2_X1 slo__sro_c137 (.ZN (slo__sro_n208), .A1 (p_0[29]), .A2 (Multiplier[29]));
OAI21_X1 slo__sro_c138 (.ZN (n_30), .A (slo__sro_n209), .B1 (slo__sro_n210), .B2 (slo__sro_n208));
XNOR2_X1 slo__sro_c139 (.ZN (slo__sro_n207), .A (p_0[29]), .B (Multiplier[29]));
XNOR2_X1 slo__sro_c140 (.ZN (p_1[29]), .A (slo__sro_n455), .B (slo__sro_n207));
INV_X1 slo__sro_c239 (.ZN (slo__sro_n336), .A (n_27));
NAND2_X1 slo__sro_c240 (.ZN (slo__sro_n335), .A1 (p_0[27]), .A2 (Multiplier[27]));
NOR2_X1 slo__sro_c241 (.ZN (slo__sro_n334), .A1 (p_0[27]), .A2 (Multiplier[27]));
OAI21_X2 slo__sro_c242 (.ZN (slo__sro_n333), .A (slo__sro_n335), .B1 (slo__sro_n334), .B2 (slo__sro_n336));
XNOR2_X1 slo__sro_c243 (.ZN (slo__sro_n332), .A (p_0[27]), .B (Multiplier[27]));
XNOR2_X1 slo__sro_c244 (.ZN (p_1[27]), .A (slo__sro_n332), .B (n_27));
NAND2_X1 slo__sro_c256 (.ZN (slo__sro_n353), .A1 (p_0[25]), .A2 (Multiplier[25]));
NOR2_X1 slo__sro_c257 (.ZN (slo__sro_n352), .A1 (p_0[25]), .A2 (Multiplier[25]));
OAI21_X2 slo__sro_c258 (.ZN (n_26), .A (slo__sro_n353), .B1 (slo__sro_n352), .B2 (slo__sro_n354));
NAND2_X1 slo__sro_c328 (.ZN (slo__sro_n458), .A1 (p_0[28]), .A2 (Multiplier[28]));
NAND2_X1 slo__sro_c329 (.ZN (slo__sro_n457), .A1 (slo__sro_n333), .A2 (Multiplier[28]));
NAND2_X1 slo__sro_c330 (.ZN (slo__sro_n456), .A1 (p_0[28]), .A2 (slo__sro_n333));
NAND3_X1 slo__sro_c331 (.ZN (slo__sro_n455), .A1 (slo__sro_n456), .A2 (slo__sro_n457), .A3 (slo__sro_n458));
XNOR2_X2 slo__sro_c332 (.ZN (slo__sro_n454), .A (slo__sro_n333), .B (Multiplier[28]));
XNOR2_X1 slo__sro_c333 (.ZN (p_1[28]), .A (slo__sro_n454), .B (p_0[28]));
OAI21_X1 slo__sro_c424 (.ZN (slo__sro_n557), .A (slo__sro_n559), .B1 (slo__sro_n560), .B2 (slo__sro_n558));
XNOR2_X1 slo__sro_c425 (.ZN (slo__sro_n556), .A (p_0[15]), .B (Multiplier[15]));
XNOR2_X1 slo__sro_c426 (.ZN (p_1[15]), .A (slo__sro_n556), .B (n_15));
NAND2_X1 slo__sro_c477 (.ZN (slo__sro_n620), .A1 (p_0[14]), .A2 (Multiplier[14]));
NOR2_X1 slo__sro_c478 (.ZN (slo__sro_n619), .A1 (p_0[14]), .A2 (Multiplier[14]));
OAI21_X1 slo__sro_c479 (.ZN (n_15), .A (slo__sro_n620), .B1 (slo__sro_n621), .B2 (slo__sro_n619));
XNOR2_X1 slo__sro_c480 (.ZN (slo__sro_n618), .A (p_0[14]), .B (Multiplier[14]));
XNOR2_X1 slo__sro_c481 (.ZN (p_1[14]), .A (slo__sro_n618), .B (n_14));
OAI21_X1 slo__sro_c498 (.ZN (slo__sro_n638), .A (p_0[26]), .B1 (n_26), .B2 (Multiplier[26]));
NAND2_X1 slo__sro_c499 (.ZN (n_27), .A1 (slo__sro_n638), .A2 (slo__sro_n639));
XNOR2_X1 slo__sro_c500 (.ZN (slo__sro_n637), .A (n_26), .B (Multiplier[26]));
XNOR2_X1 slo__sro_c501 (.ZN (p_1[26]), .A (slo__sro_n637), .B (p_0[26]));
NOR2_X1 slo__sro_c579 (.ZN (slo__sro_n744), .A1 (p_0[12]), .A2 (Multiplier[12]));
OAI21_X1 slo__sro_c580 (.ZN (slo__sro_n743), .A (slo__sro_n745), .B1 (slo__sro_n746), .B2 (slo__sro_n744));
XNOR2_X1 slo__sro_c581 (.ZN (slo__sro_n742), .A (p_0[12]), .B (Multiplier[12]));
XNOR2_X1 slo__sro_c582 (.ZN (p_1[12]), .A (slo__sro_n742), .B (n_12));
INV_X1 CLOCK_slo__sro_c1125 (.ZN (CLOCK_slo__sro_n1460), .A (slo__sro_n177));
NAND2_X1 CLOCK_slo__sro_c1126 (.ZN (CLOCK_slo__sro_n1459), .A1 (p_0[10]), .A2 (Multiplier[10]));
OAI21_X1 CLOCK_slo__sro_c1128 (.ZN (CLOCK_slo__sro_n1457), .A (CLOCK_slo__sro_n1459)
    , .B1 (CLOCK_slo__sro_n1460), .B2 (CLOCK_slo__sro_n1458));
XNOR2_X2 CLOCK_slo__sro_c1129 (.ZN (CLOCK_slo__sro_n1456), .A (p_0[10]), .B (Multiplier[10]));
XNOR2_X1 CLOCK_slo__sro_c1130 (.ZN (p_1[10]), .A (CLOCK_slo__sro_n1456), .B (slo__sro_n177));
NAND2_X1 CLOCK_slo__sro_c1143 (.ZN (CLOCK_slo__sro_n1477), .A1 (p_0[7]), .A2 (Multiplier[7]));
NOR2_X2 CLOCK_slo__sro_c1144 (.ZN (CLOCK_slo__sro_n1476), .A1 (p_0[7]), .A2 (Multiplier[7]));
OAI21_X2 CLOCK_slo__sro_c1145 (.ZN (n_8), .A (CLOCK_slo__sro_n1477), .B1 (CLOCK_slo__sro_n1478), .B2 (CLOCK_slo__sro_n1476));
XNOR2_X1 CLOCK_slo__sro_c1146 (.ZN (CLOCK_slo__sro_n1475), .A (p_0[7]), .B (Multiplier[7]));
XNOR2_X1 CLOCK_slo__sro_c1147 (.ZN (p_1[7]), .A (n_7), .B (CLOCK_slo__sro_n1475));
NAND2_X1 CLOCK_slo__sro_c1159 (.ZN (CLOCK_slo__sro_n1495), .A1 (p_0[19]), .A2 (Multiplier[19]));
INV_X2 slo__sro_c407 (.ZN (slo__sro_n546), .A (p_0[1]));
NAND2_X1 slo__sro_c408 (.ZN (slo__sro_n545), .A1 (n_1), .A2 (Multiplier[1]));
NOR2_X2 slo__sro_c409 (.ZN (slo__sro_n544), .A1 (n_1), .A2 (Multiplier[1]));
OAI21_X2 slo__sro_c410 (.ZN (n_2), .A (slo__sro_n545), .B1 (slo__sro_n546), .B2 (slo__sro_n544));
XNOR2_X1 slo__sro_c411 (.ZN (slo__sro_n543), .A (n_1), .B (Multiplier[1]));
XNOR2_X1 slo__sro_c412 (.ZN (p_1[1]), .A (slo__sro_n543), .B (p_0[1]));
OAI21_X2 CLOCK_slo__sro_c1161 (.ZN (CLOCK_slo__sro_n1493), .A (CLOCK_slo__sro_n1495)
    , .B1 (CLOCK_slo__sro_n1496), .B2 (CLOCK_slo__sro_n1494));
XNOR2_X1 CLOCK_slo__sro_c1162 (.ZN (CLOCK_slo__sro_n1492), .A (p_0[19]), .B (Multiplier[19]));
XNOR2_X1 CLOCK_slo__sro_c1163 (.ZN (p_1[19]), .A (CLOCK_slo__sro_n1492), .B (n_19));
XNOR2_X2 CLOCK_slo__mro_c1173 (.ZN (p_1[25]), .A (CLOCK_slo__mro_n1800), .B (n_25));
XNOR2_X2 CLOCK_slo__mro_c1436 (.ZN (CLOCK_slo__mro_n1800), .A (p_0[25]), .B (Multiplier[25]));

endmodule //datapath__0_116

module datapath__0_112 (p_0, p_1, p_2);

output [31:0] p_2;
input [31:0] p_0;
input [31:0] p_1;
wire CLOCK_slo__sro_n1148;
wire n_1;
wire n_2;
wire n_3;
wire n_4;
wire n_5;
wire n_6;
wire CLOCK_slo__mro_n763;
wire n_8;
wire n_9;
wire n_10;
wire n_11;
wire n_14;
wire n_15;
wire CLOCK_slo__sro_n868;
wire n_17;
wire n_18;
wire n_19;
wire n_20;
wire n_21;
wire n_22;
wire n_23;
wire n_25;
wire n_26;
wire n_27;
wire n_28;
wire n_29;
wire n_30;
wire n_32;
wire n_0;
wire n_34;
wire n_33;
wire slo__sro_n63;
wire slo__sro_n64;
wire slo__sro_n65;
wire slo__sro_n66;
wire slo__sro_n67;
wire slo__sro_n96;
wire slo__sro_n97;
wire slo__sro_n98;
wire slo__sro_n99;
wire slo__sro_n115;
wire slo__sro_n116;
wire slo__sro_n117;
wire slo__sro_n129;
wire slo__sro_n130;
wire slo__sro_n131;
wire slo__sro_n132;
wire slo__sro_n142;
wire slo__sro_n143;
wire slo__sro_n144;
wire slo__sro_n145;
wire slo__sro_n206;
wire slo__sro_n207;
wire slo__sro_n208;
wire slo__sro_n209;
wire slo__sro_n295;
wire slo__sro_n296;
wire slo__sro_n297;
wire slo__sro_n298;
wire slo__sro_n299;
wire slo__sro_n389;
wire slo__sro_n390;
wire slo__sro_n391;
wire slo__sro_n392;
wire slo__sro_n404;
wire slo__sro_n405;
wire slo__sro_n406;
wire slo__sro_n407;
wire slo__sro_n457;
wire slo__sro_n458;
wire slo__sro_n459;
wire slo__sro_n460;
wire slo__sro_n461;
wire slo__sro_n372;
wire slo__sro_n373;
wire slo__sro_n374;
wire slo__sro_n375;
wire slo__sro_n376;
wire slo__sro_n606;
wire slo__sro_n607;
wire slo__sro_n608;
wire CLOCK_slo__mro_n752;
wire CLOCK_slo__sro_n869;
wire CLOCK_slo__sro_n870;
wire CLOCK_slo__sro_n871;
wire CLOCK_slo__sro_n830;
wire CLOCK_slo__sro_n831;
wire CLOCK_slo__mro_n881;
wire CLOCK_slo__sro_n1013;
wire CLOCK_slo__sro_n1014;
wire CLOCK_slo__sro_n1015;
wire CLOCK_slo__sro_n1016;
wire CLOCK_slo__sro_n1149;
wire CLOCK_slo__sro_n1150;
wire CLOCK_slo__sro_n1151;


INV_X1 i_36 (.ZN (n_34), .A (p_0[30]));
INV_X1 i_35 (.ZN (n_33), .A (p_1[30]));
INV_X1 i_34 (.ZN (n_32), .A (n_30));
INV_X1 slo__sro_c279 (.ZN (slo__sro_n392), .A (n_10));
XOR2_X1 i_32 (.Z (p_2[31]), .A (slo__sro_n295), .B (p_0[31]));
OAI22_X1 i_31 (.ZN (n_0), .A1 (n_34), .A2 (p_1[30]), .B1 (p_0[30]), .B2 (n_33));
XNOR2_X1 i_0 (.ZN (p_2[30]), .A (n_32), .B (n_0));
FA_X1 i_30 (.CO (n_30), .S (p_2[29]), .A (p_0[29]), .B (p_1[29]), .CI (n_29));
INV_X1 slo__sro_c315 (.ZN (slo__sro_n461), .A (n_23));
FA_X1 i_28 (.CO (n_28), .S (p_2[27]), .A (p_0[27]), .B (p_1[27]), .CI (n_27));
INV_X1 CLOCK_slo__sro_c785 (.ZN (CLOCK_slo__sro_n1151), .A (n_18));
INV_X1 slo__sro_c188 (.ZN (slo__sro_n299), .A (n_30));
FA_X1 i_25 (.CO (n_25), .S (p_2[24]), .A (p_0[24]), .B (p_1[24]), .CI (slo__sro_n458));
FA_X1 i_23 (.CO (n_23), .S (p_2[22]), .A (p_0[22]), .B (p_1[22]), .CI (n_22));
FA_X1 i_22 (.CO (n_22), .S (p_2[21]), .A (p_0[21]), .B (p_1[21]), .CI (n_21));
FA_X1 i_21 (.CO (n_21), .S (p_2[20]), .A (p_0[20]), .B (p_1[20]), .CI (n_20));
FA_X1 i_20 (.CO (n_20), .S (p_2[19]), .A (p_0[19]), .B (p_1[19]), .CI (n_19));
FA_X1 i_18 (.CO (n_18), .S (p_2[17]), .A (p_0[17]), .B (p_1[17]), .CI (n_17));
FA_X1 i_17 (.CO (n_17), .S (p_2[16]), .A (p_0[16]), .B (p_1[16]), .CI (slo__sro_n64));
INV_X1 slo__sro_c28 (.ZN (slo__sro_n99), .A (n_6));
XNOR2_X1 CLOCK_slo__mro_c556 (.ZN (CLOCK_slo__mro_n881), .A (n_11), .B (p_0[11]));
FA_X1 i_14 (.CO (n_14), .S (p_2[13]), .A (p_0[13]), .B (p_1[13]), .CI (slo__sro_n373));
NOR2_X1 CLOCK_slo__sro_c787 (.ZN (CLOCK_slo__sro_n1149), .A1 (p_1[18]), .A2 (p_0[18]));
XNOR2_X2 CLOCK_slo__mro_c429 (.ZN (CLOCK_slo__mro_n752), .A (p_1[5]), .B (p_0[5]));
INV_X1 slo__sro_c293 (.ZN (slo__sro_n407), .A (n_28));
FA_X1 i_10 (.CO (n_10), .S (p_2[9]), .A (p_0[9]), .B (p_1[9]), .CI (n_9));
INV_X2 slo__sro_c72 (.ZN (slo__sro_n145), .A (n_3));
FA_X1 i_8 (.CO (n_8), .S (p_2[7]), .A (p_0[7]), .B (p_1[7]), .CI (slo__sro_n96));
INV_X1 slo__sro_c44 (.ZN (slo__sro_n117), .A (n_5));
INV_X1 slo__sro_c58 (.ZN (slo__sro_n132), .A (n_8));
FA_X1 i_5 (.CO (n_5), .S (p_2[4]), .A (p_0[4]), .B (p_1[4]), .CI (n_4));
INV_X1 slo__sro_c132 (.ZN (slo__sro_n209), .A (n_25));
FA_X1 i_3 (.CO (n_3), .S (p_2[2]), .A (p_0[2]), .B (p_1[2]), .CI (n_2));
FA_X1 i_2 (.CO (n_2), .S (p_2[1]), .A (p_0[1]), .B (p_1[1]), .CI (n_1));
XNOR2_X1 CLOCK_slo__mro_c557 (.ZN (p_2[11]), .A (CLOCK_slo__mro_n881), .B (p_1[11]));
INV_X1 slo__sro_c1 (.ZN (slo__sro_n67), .A (n_15));
NAND2_X1 slo__sro_c2 (.ZN (slo__sro_n66), .A1 (p_1[15]), .A2 (p_0[15]));
NOR2_X1 slo__sro_c3 (.ZN (slo__sro_n65), .A1 (p_1[15]), .A2 (p_0[15]));
OAI21_X1 slo__sro_c4 (.ZN (slo__sro_n64), .A (slo__sro_n66), .B1 (slo__sro_n67), .B2 (slo__sro_n65));
XNOR2_X1 slo__sro_c5 (.ZN (slo__sro_n63), .A (p_1[15]), .B (p_0[15]));
XNOR2_X1 slo__sro_c6 (.ZN (p_2[15]), .A (slo__sro_n63), .B (n_15));
NAND2_X1 slo__sro_c29 (.ZN (slo__sro_n98), .A1 (p_1[6]), .A2 (p_0[6]));
NOR2_X1 slo__sro_c30 (.ZN (slo__sro_n97), .A1 (p_1[6]), .A2 (p_0[6]));
OAI21_X1 slo__sro_c31 (.ZN (slo__sro_n96), .A (slo__sro_n98), .B1 (slo__sro_n99), .B2 (slo__sro_n97));
INV_X1 CLOCK_slo__sro_c542 (.ZN (CLOCK_slo__sro_n871), .A (n_14));
NAND2_X1 CLOCK_slo__sro_c543 (.ZN (CLOCK_slo__sro_n870), .A1 (p_1[14]), .A2 (p_0[14]));
NAND2_X1 slo__sro_c45 (.ZN (slo__sro_n116), .A1 (p_1[5]), .A2 (p_0[5]));
NOR2_X1 slo__sro_c46 (.ZN (slo__sro_n115), .A1 (p_1[5]), .A2 (p_0[5]));
OAI21_X2 slo__sro_c47 (.ZN (n_6), .A (slo__sro_n116), .B1 (slo__sro_n117), .B2 (slo__sro_n115));
XNOR2_X2 CLOCK_slo__mro_c437 (.ZN (CLOCK_slo__mro_n763), .A (n_6), .B (p_0[6]));
XNOR2_X2 CLOCK_slo__mro_c438 (.ZN (p_2[6]), .A (CLOCK_slo__mro_n763), .B (p_1[6]));
NAND2_X1 slo__sro_c59 (.ZN (slo__sro_n131), .A1 (p_1[8]), .A2 (p_0[8]));
NOR2_X1 slo__sro_c60 (.ZN (slo__sro_n130), .A1 (p_1[8]), .A2 (p_0[8]));
OAI21_X1 slo__sro_c61 (.ZN (n_9), .A (slo__sro_n131), .B1 (slo__sro_n132), .B2 (slo__sro_n130));
XNOR2_X1 slo__sro_c62 (.ZN (slo__sro_n129), .A (p_1[8]), .B (p_0[8]));
XNOR2_X1 slo__sro_c63 (.ZN (p_2[8]), .A (slo__sro_n129), .B (n_8));
NAND2_X1 slo__sro_c73 (.ZN (slo__sro_n144), .A1 (p_1[3]), .A2 (p_0[3]));
NOR2_X1 slo__sro_c74 (.ZN (slo__sro_n143), .A1 (p_1[3]), .A2 (p_0[3]));
OAI21_X2 slo__sro_c75 (.ZN (n_4), .A (slo__sro_n144), .B1 (slo__sro_n145), .B2 (slo__sro_n143));
XNOR2_X2 slo__sro_c76 (.ZN (slo__sro_n142), .A (p_1[3]), .B (p_0[3]));
XNOR2_X1 slo__sro_c77 (.ZN (p_2[3]), .A (slo__sro_n142), .B (n_3));
NAND2_X1 slo__sro_c133 (.ZN (slo__sro_n208), .A1 (p_1[25]), .A2 (p_0[25]));
NOR2_X1 slo__sro_c134 (.ZN (slo__sro_n207), .A1 (p_1[25]), .A2 (p_0[25]));
OAI21_X1 slo__sro_c135 (.ZN (n_26), .A (slo__sro_n208), .B1 (slo__sro_n209), .B2 (slo__sro_n207));
XNOR2_X1 slo__sro_c136 (.ZN (slo__sro_n206), .A (p_1[25]), .B (p_0[25]));
XNOR2_X1 slo__sro_c137 (.ZN (p_2[25]), .A (slo__sro_n206), .B (n_25));
NOR2_X1 slo__sro_c189 (.ZN (slo__sro_n298), .A1 (n_33), .A2 (p_0[30]));
NAND2_X1 slo__sro_c190 (.ZN (slo__sro_n297), .A1 (slo__sro_n298), .A2 (slo__sro_n299));
OR2_X1 slo__sro_c191 (.ZN (slo__sro_n296), .A1 (p_1[30]), .A2 (n_34));
OAI21_X1 slo__sro_c192 (.ZN (slo__sro_n295), .A (slo__sro_n297), .B1 (n_32), .B2 (slo__sro_n296));
NAND2_X1 slo__sro_c280 (.ZN (slo__sro_n391), .A1 (p_1[10]), .A2 (p_0[10]));
NOR2_X1 slo__sro_c281 (.ZN (slo__sro_n390), .A1 (p_1[10]), .A2 (p_0[10]));
OAI21_X1 CLOCK_slo__sro_c730 (.ZN (slo__sro_n607), .A (n_11), .B1 (p_1[11]), .B2 (p_0[11]));
XNOR2_X1 slo__sro_c283 (.ZN (slo__sro_n389), .A (p_1[10]), .B (p_0[10]));
XNOR2_X1 slo__sro_c284 (.ZN (p_2[10]), .A (slo__sro_n389), .B (n_10));
NAND2_X1 slo__sro_c294 (.ZN (slo__sro_n406), .A1 (p_1[28]), .A2 (p_0[28]));
NOR2_X1 slo__sro_c295 (.ZN (slo__sro_n405), .A1 (p_1[28]), .A2 (p_0[28]));
OAI21_X1 slo__sro_c296 (.ZN (n_29), .A (slo__sro_n406), .B1 (slo__sro_n407), .B2 (slo__sro_n405));
XNOR2_X1 slo__sro_c297 (.ZN (slo__sro_n404), .A (p_1[28]), .B (p_0[28]));
XNOR2_X2 slo__sro_c298 (.ZN (p_2[28]), .A (slo__sro_n404), .B (n_28));
NAND2_X1 slo__sro_c316 (.ZN (slo__sro_n460), .A1 (p_1[23]), .A2 (p_0[23]));
NOR2_X1 slo__sro_c317 (.ZN (slo__sro_n459), .A1 (p_1[23]), .A2 (p_0[23]));
OAI21_X1 slo__sro_c318 (.ZN (slo__sro_n458), .A (slo__sro_n460), .B1 (slo__sro_n461), .B2 (slo__sro_n459));
XNOR2_X1 slo__sro_c319 (.ZN (slo__sro_n457), .A (p_1[23]), .B (p_0[23]));
XNOR2_X1 slo__sro_c320 (.ZN (p_2[23]), .A (slo__sro_n457), .B (n_23));
NAND2_X1 slo__sro_c387 (.ZN (slo__sro_n608), .A1 (p_1[11]), .A2 (p_0[11]));
INV_X1 slo__sro_c265 (.ZN (slo__sro_n376), .A (slo__sro_n606));
NAND2_X1 slo__sro_c266 (.ZN (slo__sro_n375), .A1 (p_1[12]), .A2 (p_0[12]));
NOR2_X1 slo__sro_c267 (.ZN (slo__sro_n374), .A1 (p_1[12]), .A2 (p_0[12]));
OAI21_X1 slo__sro_c268 (.ZN (slo__sro_n373), .A (slo__sro_n375), .B1 (slo__sro_n376), .B2 (slo__sro_n374));
XNOR2_X1 slo__sro_c269 (.ZN (slo__sro_n372), .A (p_1[12]), .B (p_0[12]));
XNOR2_X1 slo__sro_c270 (.ZN (p_2[12]), .A (slo__sro_n372), .B (slo__sro_n606));
NAND2_X1 slo__sro_c389 (.ZN (slo__sro_n606), .A1 (slo__sro_n607), .A2 (slo__sro_n608));
OAI21_X2 CLOCK_slo__sro_c720 (.ZN (n_11), .A (slo__sro_n391), .B1 (slo__sro_n392), .B2 (slo__sro_n390));
INV_X1 CLOCK_slo__sro_c645 (.ZN (CLOCK_slo__sro_n1016), .A (p_1[26]));
XNOR2_X1 CLOCK_slo__mro_c430 (.ZN (p_2[5]), .A (CLOCK_slo__mro_n752), .B (n_5));
NOR2_X1 CLOCK_slo__sro_c544 (.ZN (CLOCK_slo__sro_n869), .A1 (p_1[14]), .A2 (p_0[14]));
OAI21_X1 CLOCK_slo__sro_c545 (.ZN (n_15), .A (CLOCK_slo__sro_n870), .B1 (CLOCK_slo__sro_n871), .B2 (CLOCK_slo__sro_n869));
XNOR2_X1 CLOCK_slo__sro_c546 (.ZN (CLOCK_slo__sro_n868), .A (p_1[14]), .B (p_0[14]));
XNOR2_X1 CLOCK_slo__sro_c547 (.ZN (p_2[14]), .A (CLOCK_slo__sro_n868), .B (n_14));
INV_X1 CLOCK_slo__sro_c503 (.ZN (CLOCK_slo__sro_n831), .A (p_0[0]));
INV_X2 CLOCK_slo__sro_c504 (.ZN (CLOCK_slo__sro_n830), .A (p_1[0]));
NOR2_X2 CLOCK_slo__sro_c505 (.ZN (n_1), .A1 (CLOCK_slo__sro_n830), .A2 (CLOCK_slo__sro_n831));
XNOR2_X1 CLOCK_slo__sro_c506 (.ZN (p_2[0]), .A (p_1[0]), .B (CLOCK_slo__sro_n831));
NAND2_X1 CLOCK_slo__sro_c646 (.ZN (CLOCK_slo__sro_n1015), .A1 (n_26), .A2 (p_0[26]));
NOR2_X1 CLOCK_slo__sro_c647 (.ZN (CLOCK_slo__sro_n1014), .A1 (n_26), .A2 (p_0[26]));
OAI21_X1 CLOCK_slo__sro_c648 (.ZN (n_27), .A (CLOCK_slo__sro_n1015), .B1 (CLOCK_slo__sro_n1016), .B2 (CLOCK_slo__sro_n1014));
XNOR2_X1 CLOCK_slo__sro_c649 (.ZN (CLOCK_slo__sro_n1013), .A (n_26), .B (p_0[26]));
XNOR2_X1 CLOCK_slo__sro_c650 (.ZN (p_2[26]), .A (CLOCK_slo__sro_n1013), .B (p_1[26]));
NAND2_X1 CLOCK_slo__sro_c786 (.ZN (CLOCK_slo__sro_n1150), .A1 (p_1[18]), .A2 (p_0[18]));
OAI21_X1 CLOCK_slo__sro_c788 (.ZN (n_19), .A (CLOCK_slo__sro_n1150), .B1 (CLOCK_slo__sro_n1151), .B2 (CLOCK_slo__sro_n1149));
XNOR2_X1 CLOCK_slo__sro_c789 (.ZN (CLOCK_slo__sro_n1148), .A (p_1[18]), .B (p_0[18]));
XNOR2_X1 CLOCK_slo__sro_c790 (.ZN (p_2[18]), .A (CLOCK_slo__sro_n1148), .B (n_18));

endmodule //datapath__0_112

module datapath__0_111 (p_0_17_PP_0, Multiplier, p_0, p_1);

output [31:0] p_1;
input [31:0] Multiplier;
input [31:0] p_0;
input p_0_17_PP_0;
wire slo__sro_n339;
wire slo__sro_n338;
wire n_2;
wire n_3;
wire n_4;
wire n_5;
wire n_6;
wire n_8;
wire n_9;
wire n_10;
wire n_11;
wire n_14;
wire n_15;
wire n_16;
wire n_19;
wire n_20;
wire n_21;
wire CLOCK_slo__sro_n1148;
wire n_23;
wire n_25;
wire n_26;
wire n_27;
wire n_28;
wire n_29;
wire n_30;
wire n_32;
wire n_0;
wire n_34;
wire n_33;
wire n_31;
wire slo__sro_n185;
wire slo__sro_n186;
wire slo__sro_n187;
wire slo__sro_n188;
wire slo__sro_n189;
wire slo__sro_n202;
wire slo__sro_n203;
wire slo__sro_n204;
wire slo__sro_n205;
wire slo__sro_n217;
wire slo__sro_n218;
wire slo__sro_n219;
wire slo__sro_n220;
wire slo__sro_n221;
wire slo__sro_n672;
wire slo__sro_n298;
wire slo__sro_n299;
wire slo__sro_n300;
wire slo__sro_n301;
wire slo__sro_n314;
wire slo__sro_n315;
wire slo__sro_n316;
wire slo__sro_n317;
wire slo__sro_n340;
wire slo__sro_n341;
wire slo__mro_n630;
wire slo__sro_n673;
wire slo__sro_n674;
wire slo__sro_n675;
wire slo__sro_n676;
wire slo__sro_n945;
wire slo__sro_n946;
wire slo__sro_n947;
wire CLOCK_slo__sro_n1122;
wire CLOCK_slo__sro_n1123;
wire CLOCK_slo__sro_n1124;
wire CLOCK_slo__sro_n1125;
wire CLOCK_slo__sro_n1126;
wire CLOCK_slo__sro_n1146;
wire CLOCK_slo__sro_n1147;
wire slo__sro_n457;
wire slo__sro_n458;
wire slo__sro_n459;
wire slo__sro_n460;
wire slo__sro_n461;
wire slo__sro_n563;
wire slo__sro_n564;
wire slo__sro_n565;
wire slo__sro_n566;
wire slo__sro_n567;
wire CLOCK_slo__sro_n1149;
wire CLOCK_slo__sro_n1150;
wire CLOCK_slo__sro_n1214;
wire CLOCK_slo__sro_n1215;
wire CLOCK_slo__sro_n1216;
wire CLOCK_slo__sro_n1217;
wire CLOCK_slo__sro_n1246;
wire CLOCK_slo__sro_n1247;
wire CLOCK_slo__sro_n1248;
wire CLOCK_slo__sro_n1249;
wire CLOCK_slo__sro_n1393;
wire CLOCK_slo__sro_n1394;
wire CLOCK_slo__sro_n1395;
wire CLOCK_slo__sro_n1396;


INV_X1 i_36 (.ZN (n_34), .A (Multiplier[30]));
INV_X1 i_35 (.ZN (n_33), .A (p_0[30]));
INV_X1 i_34 (.ZN (n_32), .A (n_30));
XNOR2_X2 slo__mro_c501 (.ZN (slo__mro_n630), .A (n_23), .B (Multiplier[23]));
XOR2_X1 i_32 (.Z (p_1[31]), .A (Multiplier[31]), .B (n_31));
OAI22_X1 i_31 (.ZN (n_0), .A1 (n_34), .A2 (p_0[30]), .B1 (n_33), .B2 (Multiplier[30]));
XNOR2_X1 i_0 (.ZN (p_1[30]), .A (n_32), .B (n_0));
NAND2_X1 slo__sro_c218 (.ZN (slo__sro_n316), .A1 (p_0[23]), .A2 (Multiplier[23]));
INV_X1 CLOCK_slo__sro_c995 (.ZN (CLOCK_slo__sro_n1249), .A (n_5));
FA_X1 i_28 (.CO (n_28), .S (p_1[27]), .A (Multiplier[27]), .B (p_0[27]), .CI (n_27));
FA_X1 i_27 (.CO (n_27), .S (p_1[26]), .A (Multiplier[26]), .B (p_0[26]), .CI (n_26));
FA_X1 i_26 (.CO (n_26), .S (p_1[25]), .A (Multiplier[25]), .B (p_0[25]), .CI (n_25));
FA_X1 i_25 (.CO (n_25), .S (p_1[24]), .A (Multiplier[24]), .B (p_0[24]), .CI (slo__sro_n314));
NOR2_X1 slo__sro_c236 (.ZN (slo__sro_n340), .A1 (n_33), .A2 (Multiplier[30]));
INV_X1 slo__sro_c764 (.ZN (slo__sro_n947), .A (Multiplier[0]));
XNOR2_X1 CLOCK_slo__sro_c910 (.ZN (CLOCK_slo__sro_n1146), .A (p_0[16]), .B (Multiplier[16]));
FA_X1 i_21 (.CO (n_21), .S (p_1[20]), .A (Multiplier[20]), .B (p_0[20]), .CI (n_20));
FA_X1 i_20 (.CO (n_20), .S (p_1[19]), .A (Multiplier[19]), .B (p_0[19]), .CI (n_19));
INV_X1 slo__sro_c134 (.ZN (slo__sro_n205), .A (slo__sro_n218));
NAND2_X1 CLOCK_slo__sro_c1100 (.ZN (CLOCK_slo__sro_n1395), .A1 (p_0[18]), .A2 (Multiplier[18]));
FA_X1 i_16 (.CO (n_16), .S (p_1[15]), .A (Multiplier[15]), .B (p_0[15]), .CI (n_15));
FA_X1 i_15 (.CO (n_15), .S (p_1[14]), .A (Multiplier[14]), .B (p_0[14]), .CI (n_14));
FA_X1 i_14 (.CO (n_14), .S (p_1[13]), .A (Multiplier[13]), .B (p_0[13]), .CI (slo__sro_n458));
OAI21_X2 CLOCK_slo__sro_c909 (.ZN (CLOCK_slo__sro_n1147), .A (CLOCK_slo__sro_n1149)
    , .B1 (CLOCK_slo__sro_n1150), .B2 (CLOCK_slo__sro_n1148));
INV_X1 CLOCK_slo__sro_c906 (.ZN (CLOCK_slo__sro_n1150), .A (n_16));
FA_X1 i_11 (.CO (n_11), .S (p_1[10]), .A (Multiplier[10]), .B (p_0[10]), .CI (n_10));
FA_X1 i_10 (.CO (n_10), .S (p_1[9]), .A (Multiplier[9]), .B (p_0[9]), .CI (n_9));
FA_X1 i_9 (.CO (n_9), .S (p_1[8]), .A (Multiplier[8]), .B (p_0[8]), .CI (n_8));
INV_X1 slo__sro_c150 (.ZN (slo__sro_n221), .A (n_6));
INV_X1 slo__sro_c235 (.ZN (slo__sro_n341), .A (n_30));
FA_X1 i_5 (.CO (n_5), .S (p_1[4]), .A (Multiplier[4]), .B (p_0[4]), .CI (n_4));
FA_X1 i_4 (.CO (n_4), .S (p_1[3]), .A (Multiplier[3]), .B (p_0[3]), .CI (n_3));
FA_X1 i_3 (.CO (n_3), .S (p_1[2]), .A (Multiplier[2]), .B (p_0[2]), .CI (n_2));
FA_X1 i_2 (.CO (n_2), .S (p_1[1]), .A (Multiplier[1]), .B (p_0[1]), .CI (slo__sro_n945));
INV_X1 CLOCK_slo__sro_c882 (.ZN (CLOCK_slo__sro_n1126), .A (n_11));
INV_X2 slo__sro_c120 (.ZN (slo__sro_n189), .A (CLOCK_slo__sro_n1147));
NAND2_X1 slo__sro_c121 (.ZN (slo__sro_n188), .A1 (p_0[17]), .A2 (Multiplier[17]));
NOR2_X1 slo__sro_c122 (.ZN (slo__sro_n187), .A1 (p_0[17]), .A2 (Multiplier[17]));
OAI21_X1 slo__sro_c123 (.ZN (slo__sro_n186), .A (slo__sro_n188), .B1 (slo__sro_n189), .B2 (slo__sro_n187));
XNOR2_X1 slo__sro_c124 (.ZN (slo__sro_n185), .A (p_0_17_PP_0), .B (Multiplier[17]));
XNOR2_X1 slo__sro_c125 (.ZN (p_1[17]), .A (slo__sro_n185), .B (CLOCK_slo__sro_n1147));
NAND2_X1 slo__sro_c135 (.ZN (slo__sro_n204), .A1 (p_0[7]), .A2 (Multiplier[7]));
NOR2_X1 slo__sro_c136 (.ZN (slo__sro_n203), .A1 (p_0[7]), .A2 (Multiplier[7]));
OAI21_X1 slo__sro_c137 (.ZN (n_8), .A (slo__sro_n204), .B1 (slo__sro_n205), .B2 (slo__sro_n203));
XNOR2_X2 slo__sro_c138 (.ZN (slo__sro_n202), .A (p_0[7]), .B (Multiplier[7]));
XNOR2_X2 slo__sro_c139 (.ZN (p_1[7]), .A (slo__sro_n202), .B (slo__sro_n218));
NAND2_X1 slo__sro_c151 (.ZN (slo__sro_n220), .A1 (p_0[6]), .A2 (Multiplier[6]));
NOR2_X1 slo__sro_c152 (.ZN (slo__sro_n219), .A1 (p_0[6]), .A2 (Multiplier[6]));
OAI21_X2 slo__sro_c153 (.ZN (slo__sro_n218), .A (slo__sro_n220), .B1 (slo__sro_n221), .B2 (slo__sro_n219));
XNOR2_X1 slo__sro_c154 (.ZN (slo__sro_n217), .A (p_0[6]), .B (Multiplier[6]));
XNOR2_X1 slo__sro_c155 (.ZN (p_1[6]), .A (slo__sro_n217), .B (n_6));
INV_X1 slo__sro_c217 (.ZN (slo__sro_n317), .A (n_23));
INV_X1 slo__sro_c201 (.ZN (slo__sro_n301), .A (n_29));
NAND2_X1 slo__sro_c202 (.ZN (slo__sro_n300), .A1 (p_0[29]), .A2 (Multiplier[29]));
NOR2_X1 slo__sro_c203 (.ZN (slo__sro_n299), .A1 (p_0[29]), .A2 (Multiplier[29]));
OAI21_X1 slo__sro_c204 (.ZN (n_30), .A (slo__sro_n300), .B1 (slo__sro_n301), .B2 (slo__sro_n299));
XNOR2_X1 slo__sro_c205 (.ZN (slo__sro_n298), .A (p_0[29]), .B (Multiplier[29]));
XNOR2_X1 slo__sro_c206 (.ZN (p_1[29]), .A (n_29), .B (slo__sro_n298));
NOR2_X1 slo__sro_c219 (.ZN (slo__sro_n315), .A1 (p_0[23]), .A2 (Multiplier[23]));
OAI21_X1 slo__sro_c220 (.ZN (slo__sro_n314), .A (slo__sro_n316), .B1 (slo__sro_n317), .B2 (slo__sro_n315));
BUF_X2 slo__sro_c539 (.Z (slo__sro_n676), .A (slo__sro_n564));
NAND2_X1 slo__sro_c540 (.ZN (slo__sro_n675), .A1 (p_0[22]), .A2 (Multiplier[22]));
NAND2_X1 slo__sro_c237 (.ZN (slo__sro_n339), .A1 (slo__sro_n340), .A2 (slo__sro_n341));
OR2_X1 slo__sro_c238 (.ZN (slo__sro_n338), .A1 (p_0[30]), .A2 (n_34));
OAI21_X1 slo__sro_c239 (.ZN (n_31), .A (slo__sro_n339), .B1 (n_32), .B2 (slo__sro_n338));
XNOR2_X2 slo__mro_c502 (.ZN (p_1[23]), .A (slo__mro_n630), .B (p_0[23]));
NAND2_X4 slo__sro_c541 (.ZN (slo__sro_n674), .A1 (slo__sro_n676), .A2 (Multiplier[22]));
NAND2_X1 slo__sro_c542 (.ZN (slo__sro_n673), .A1 (slo__sro_n676), .A2 (p_0[22]));
NAND3_X2 slo__sro_c543 (.ZN (n_23), .A1 (slo__sro_n673), .A2 (slo__sro_n674), .A3 (slo__sro_n675));
XNOR2_X1 slo__sro_c544 (.ZN (slo__sro_n672), .A (p_0[22]), .B (Multiplier[22]));
XNOR2_X1 slo__sro_c545 (.ZN (p_1[22]), .A (slo__sro_n672), .B (slo__sro_n676));
INV_X2 slo__sro_c765 (.ZN (slo__sro_n946), .A (p_0[0]));
NOR2_X1 slo__sro_c766 (.ZN (slo__sro_n945), .A1 (slo__sro_n946), .A2 (slo__sro_n947));
XNOR2_X1 slo__sro_c767 (.ZN (p_1[0]), .A (p_0[0]), .B (slo__sro_n947));
NAND2_X1 CLOCK_slo__sro_c883 (.ZN (CLOCK_slo__sro_n1125), .A1 (p_0[11]), .A2 (Multiplier[11]));
NOR2_X1 CLOCK_slo__sro_c884 (.ZN (CLOCK_slo__sro_n1124), .A1 (p_0[11]), .A2 (Multiplier[11]));
OAI21_X2 CLOCK_slo__sro_c885 (.ZN (CLOCK_slo__sro_n1123), .A (CLOCK_slo__sro_n1125)
    , .B1 (CLOCK_slo__sro_n1126), .B2 (CLOCK_slo__sro_n1124));
XNOR2_X1 CLOCK_slo__sro_c886 (.ZN (CLOCK_slo__sro_n1122), .A (p_0[11]), .B (Multiplier[11]));
XNOR2_X1 CLOCK_slo__sro_c887 (.ZN (p_1[11]), .A (CLOCK_slo__sro_n1122), .B (n_11));
NAND2_X1 CLOCK_slo__sro_c907 (.ZN (CLOCK_slo__sro_n1149), .A1 (p_0[16]), .A2 (Multiplier[16]));
NOR2_X1 CLOCK_slo__sro_c908 (.ZN (CLOCK_slo__sro_n1148), .A1 (p_0[16]), .A2 (Multiplier[16]));
INV_X1 slo__sro_c351 (.ZN (slo__sro_n461), .A (CLOCK_slo__sro_n1123));
NAND2_X1 slo__sro_c352 (.ZN (slo__sro_n460), .A1 (p_0[12]), .A2 (Multiplier[12]));
NOR2_X1 slo__sro_c353 (.ZN (slo__sro_n459), .A1 (p_0[12]), .A2 (Multiplier[12]));
OAI21_X1 slo__sro_c354 (.ZN (slo__sro_n458), .A (slo__sro_n460), .B1 (slo__sro_n461), .B2 (slo__sro_n459));
XNOR2_X1 slo__sro_c355 (.ZN (slo__sro_n457), .A (p_0[12]), .B (Multiplier[12]));
XNOR2_X1 slo__sro_c356 (.ZN (p_1[12]), .A (slo__sro_n457), .B (CLOCK_slo__sro_n1123));
INV_X1 slo__sro_c449 (.ZN (slo__sro_n567), .A (n_21));
NAND2_X1 slo__sro_c450 (.ZN (slo__sro_n566), .A1 (p_0[21]), .A2 (Multiplier[21]));
NOR2_X1 slo__sro_c451 (.ZN (slo__sro_n565), .A1 (p_0[21]), .A2 (Multiplier[21]));
OAI21_X1 slo__sro_c452 (.ZN (slo__sro_n564), .A (slo__sro_n566), .B1 (slo__sro_n567), .B2 (slo__sro_n565));
XNOR2_X1 slo__sro_c453 (.ZN (slo__sro_n563), .A (p_0[21]), .B (Multiplier[21]));
XNOR2_X1 slo__sro_c454 (.ZN (p_1[21]), .A (slo__sro_n563), .B (n_21));
XNOR2_X1 CLOCK_slo__sro_c911 (.ZN (p_1[16]), .A (n_16), .B (CLOCK_slo__sro_n1146));
INV_X1 CLOCK_slo__sro_c969 (.ZN (CLOCK_slo__sro_n1217), .A (n_28));
NAND2_X1 CLOCK_slo__sro_c970 (.ZN (CLOCK_slo__sro_n1216), .A1 (p_0[28]), .A2 (Multiplier[28]));
NOR2_X1 CLOCK_slo__sro_c971 (.ZN (CLOCK_slo__sro_n1215), .A1 (p_0[28]), .A2 (Multiplier[28]));
OAI21_X2 CLOCK_slo__sro_c972 (.ZN (n_29), .A (CLOCK_slo__sro_n1216), .B1 (CLOCK_slo__sro_n1217), .B2 (CLOCK_slo__sro_n1215));
XNOR2_X1 CLOCK_slo__sro_c973 (.ZN (CLOCK_slo__sro_n1214), .A (p_0[28]), .B (Multiplier[28]));
XNOR2_X1 CLOCK_slo__sro_c974 (.ZN (p_1[28]), .A (CLOCK_slo__sro_n1214), .B (n_28));
NAND2_X1 CLOCK_slo__sro_c996 (.ZN (CLOCK_slo__sro_n1248), .A1 (p_0[5]), .A2 (Multiplier[5]));
NOR2_X1 CLOCK_slo__sro_c997 (.ZN (CLOCK_slo__sro_n1247), .A1 (p_0[5]), .A2 (Multiplier[5]));
OAI21_X2 CLOCK_slo__sro_c998 (.ZN (n_6), .A (CLOCK_slo__sro_n1248), .B1 (CLOCK_slo__sro_n1247), .B2 (CLOCK_slo__sro_n1249));
XNOR2_X1 CLOCK_slo__sro_c999 (.ZN (CLOCK_slo__sro_n1246), .A (p_0[5]), .B (Multiplier[5]));
XNOR2_X1 CLOCK_slo__sro_c1000 (.ZN (p_1[5]), .A (CLOCK_slo__sro_n1246), .B (n_5));
INV_X1 CLOCK_slo__sro_c1099 (.ZN (CLOCK_slo__sro_n1396), .A (slo__sro_n186));
NOR2_X1 CLOCK_slo__sro_c1101 (.ZN (CLOCK_slo__sro_n1394), .A1 (p_0[18]), .A2 (Multiplier[18]));
OAI21_X1 CLOCK_slo__sro_c1102 (.ZN (n_19), .A (CLOCK_slo__sro_n1395), .B1 (CLOCK_slo__sro_n1394), .B2 (CLOCK_slo__sro_n1396));
XNOR2_X1 CLOCK_slo__sro_c1103 (.ZN (CLOCK_slo__sro_n1393), .A (p_0[18]), .B (Multiplier[18]));
XNOR2_X1 CLOCK_slo__sro_c1104 (.ZN (p_1[18]), .A (CLOCK_slo__sro_n1393), .B (slo__sro_n186));

endmodule //datapath__0_111

module datapath__0_107 (p_0_9_PP_0, p_0, p_1, p_2);

output [31:0] p_2;
input [31:0] p_0;
input [31:0] p_1;
input p_0_9_PP_0;
wire CLOCK_slo__sro_n917;
wire slo__sro_n511;
wire slo__sro_n470;
wire n_1;
wire n_3;
wire n_4;
wire n_5;
wire n_6;
wire n_7;
wire n_8;
wire n_9;
wire n_10;
wire n_12;
wire n_14;
wire n_15;
wire n_19;
wire n_20;
wire n_21;
wire n_23;
wire n_25;
wire n_27;
wire n_28;
wire n_29;
wire n_30;
wire n_32;
wire n_0;
wire n_34;
wire n_33;
wire n_31;
wire slo__sro_n81;
wire slo__sro_n82;
wire slo__sro_n83;
wire slo__sro_n84;
wire slo__sro_n85;
wire slo__sro_n113;
wire slo__sro_n114;
wire slo__sro_n115;
wire slo__sro_n116;
wire slo__sro_n117;
wire slo__sro_n131;
wire slo__sro_n132;
wire slo__sro_n133;
wire slo__sro_n134;
wire slo__sro_n149;
wire slo__sro_n150;
wire slo__sro_n151;
wire slo__sro_n152;
wire slo__sro_n181;
wire slo__sro_n182;
wire slo__sro_n183;
wire slo__sro_n184;
wire slo__sro_n194;
wire slo__sro_n195;
wire slo__sro_n196;
wire slo__sro_n197;
wire slo__sro_n291;
wire slo__sro_n292;
wire slo__sro_n293;
wire slo__sro_n294;
wire slo__sro_n303;
wire slo__sro_n304;
wire slo__sro_n305;
wire slo__sro_n306;
wire slo__sro_n318;
wire slo__sro_n319;
wire slo__sro_n320;
wire slo__sro_n331;
wire slo__sro_n332;
wire slo__sro_n333;
wire slo__sro_n344;
wire slo__sro_n345;
wire slo__sro_n346;
wire slo__sro_n347;
wire slo__sro_n434;
wire slo__sro_n435;
wire slo__sro_n436;
wire slo__sro_n437;
wire slo__sro_n438;
wire slo__mro_n453;
wire slo__sro_n471;
wire slo__sro_n472;
wire slo__sro_n473;
wire slo__sro_n510;
wire slo__sro_n491;
wire slo__sro_n492;
wire slo__sro_n493;
wire slo__sro_n494;
wire slo__sro_n512;
wire slo__sro_n513;
wire CLOCK_slo__sro_n767;
wire CLOCK_slo__sro_n768;
wire CLOCK_slo__sro_n786;
wire CLOCK_slo__sro_n787;
wire CLOCK_slo__sro_n788;
wire CLOCK_slo__sro_n789;
wire CLOCK_slo__sro_n790;
wire CLOCK_slo__sro_n898;
wire CLOCK_slo__sro_n918;
wire CLOCK_slo__sro_n919;
wire CLOCK_slo__sro_n960;
wire CLOCK_slo__sro_n961;
wire CLOCK_slo__sro_n962;
wire CLOCK_slo__sro_n963;
wire CLOCK_slo__sro_n1101;
wire CLOCK_slo__sro_n1102;
wire CLOCK_slo__sro_n1103;
wire CLOCK_slo__sro_n1104;
wire CLOCK_slo__sro_n1105;


INV_X1 i_36 (.ZN (n_34), .A (p_0[30]));
INV_X1 i_35 (.ZN (n_33), .A (p_1[30]));
INV_X1 i_34 (.ZN (n_32), .A (n_30));
NAND2_X1 slo__sro_c200 (.ZN (slo__sro_n306), .A1 (p_1[21]), .A2 (p_0[21]));
INV_X1 CLOCK_slo__sro_c652 (.ZN (CLOCK_slo__sro_n919), .A (p_1[17]));
OAI22_X1 i_31 (.ZN (n_0), .A1 (n_34), .A2 (p_1[30]), .B1 (p_0[30]), .B2 (n_33));
XNOR2_X1 i_0 (.ZN (p_2[30]), .A (n_32), .B (n_0));
FA_X1 i_30 (.CO (n_30), .S (p_2[29]), .A (p_0[29]), .B (p_1[29]), .CI (n_29));
FA_X1 i_29 (.CO (n_29), .S (p_2[28]), .A (p_0[28]), .B (p_1[28]), .CI (n_28));
FA_X1 i_28 (.CO (n_28), .S (p_2[27]), .A (p_0[27]), .B (p_1[27]), .CI (n_27));
FA_X1 i_27 (.CO (n_27), .S (p_2[26]), .A (p_0[26]), .B (p_1[26]), .CI (slo__sro_n345));
XNOR2_X2 slo__mro_c316 (.ZN (slo__mro_n453), .A (n_1), .B (p_0[1]));
NAND2_X1 slo__sro_c236 (.ZN (slo__sro_n347), .A1 (p_1[25]), .A2 (p_0[25]));
NAND2_X1 slo__sro_c212 (.ZN (slo__sro_n320), .A1 (p_1[20]), .A2 (p_0[20]));
NAND2_X1 slo__sro_c224 (.ZN (slo__sro_n333), .A1 (p_1[22]), .A2 (p_0[22]));
FA_X1 i_20 (.CO (n_20), .S (p_2[19]), .A (p_0[19]), .B (p_1[19]), .CI (n_19));
FA_X1 i_19 (.CO (n_19), .S (p_2[18]), .A (p_0[18]), .B (p_1[18]), .CI (slo__sro_n492));
OAI21_X2 slo__sro_c366 (.ZN (n_3), .A (slo__sro_n512), .B1 (slo__sro_n513), .B2 (slo__sro_n511));
INV_X1 slo__sro_c58 (.ZN (slo__sro_n134), .A (n_1));
FA_X1 i_15 (.CO (n_15), .S (p_2[14]), .A (p_0[14]), .B (p_1[14]), .CI (n_14));
FA_X1 i_14 (.CO (n_14), .S (p_2[13]), .A (p_0[13]), .B (p_1[13]), .CI (CLOCK_slo__sro_n1102));
FA_X1 i_12 (.CO (n_12), .S (p_2[11]), .A (p_0[11]), .B (p_1[11]), .CI (slo__sro_n82));
INV_X1 slo__sro_c44 (.ZN (slo__sro_n117), .A (CLOCK_slo__sro_n787));
INV_X1 slo__sro_c103 (.ZN (slo__sro_n184), .A (n_7));
FA_X1 i_9 (.CO (n_9), .S (p_2[8]), .A (p_0[8]), .B (p_1[8]), .CI (n_8));
INV_X1 slo__sro_c117 (.ZN (slo__sro_n197), .A (n_4));
FA_X1 i_7 (.CO (n_7), .S (p_2[6]), .A (p_0[6]), .B (p_1[6]), .CI (n_6));
FA_X1 i_6 (.CO (n_6), .S (p_2[5]), .A (p_0[5]), .B (p_1[5]), .CI (n_5));
INV_X1 slo__sro_c188 (.ZN (slo__sro_n294), .A (n_30));
INV_X1 slo__sro_c363 (.ZN (slo__sro_n513), .A (slo__sro_n131));
INV_X1 CLOCK_slo__sro_c529 (.ZN (CLOCK_slo__sro_n768), .A (p_0[0]));
INV_X1 slo__sro_c74 (.ZN (slo__sro_n152), .A (n_9));
INV_X1 CLOCK_slo__sro_c550 (.ZN (CLOCK_slo__sro_n790), .A (n_15));
INV_X1 slo__sro_c17 (.ZN (slo__sro_n85), .A (n_10));
NAND2_X1 slo__sro_c18 (.ZN (slo__sro_n84), .A1 (p_1[10]), .A2 (p_0[10]));
NOR2_X1 slo__sro_c19 (.ZN (slo__sro_n83), .A1 (p_1[10]), .A2 (p_0[10]));
OAI21_X1 slo__sro_c20 (.ZN (slo__sro_n82), .A (slo__sro_n84), .B1 (slo__sro_n85), .B2 (slo__sro_n83));
XNOR2_X1 slo__sro_c21 (.ZN (slo__sro_n81), .A (p_1[10]), .B (p_0[10]));
XNOR2_X1 slo__sro_c22 (.ZN (p_2[10]), .A (slo__sro_n81), .B (n_10));
NAND2_X1 slo__sro_c45 (.ZN (slo__sro_n116), .A1 (p_1[16]), .A2 (p_0[16]));
NOR2_X1 slo__sro_c46 (.ZN (slo__sro_n115), .A1 (p_1[16]), .A2 (p_0[16]));
OAI21_X1 slo__sro_c47 (.ZN (slo__sro_n114), .A (slo__sro_n116), .B1 (slo__sro_n117), .B2 (slo__sro_n115));
XNOR2_X1 slo__sro_c48 (.ZN (slo__sro_n113), .A (p_1[16]), .B (p_0[16]));
XNOR2_X1 slo__sro_c49 (.ZN (p_2[16]), .A (slo__sro_n113), .B (CLOCK_slo__sro_n787));
NAND2_X1 slo__sro_c59 (.ZN (slo__sro_n133), .A1 (p_1[1]), .A2 (p_0[1]));
NOR2_X1 slo__sro_c60 (.ZN (slo__sro_n132), .A1 (p_1[1]), .A2 (p_0[1]));
OAI21_X2 slo__sro_c61 (.ZN (slo__sro_n131), .A (slo__sro_n133), .B1 (slo__sro_n132), .B2 (slo__sro_n134));
INV_X2 slo__sro_c326 (.ZN (slo__sro_n473), .A (n_3));
NAND2_X1 slo__sro_c327 (.ZN (slo__sro_n472), .A1 (p_1[3]), .A2 (p_0[3]));
NAND2_X1 slo__sro_c75 (.ZN (slo__sro_n151), .A1 (p_1[9]), .A2 (p_0_9_PP_0));
NOR2_X1 slo__sro_c76 (.ZN (slo__sro_n150), .A1 (p_1[9]), .A2 (p_0[9]));
OAI21_X1 slo__sro_c77 (.ZN (n_10), .A (slo__sro_n151), .B1 (slo__sro_n152), .B2 (slo__sro_n150));
XNOR2_X1 slo__sro_c78 (.ZN (slo__sro_n149), .A (p_1[9]), .B (p_0[9]));
XNOR2_X1 slo__sro_c79 (.ZN (p_2[9]), .A (slo__sro_n149), .B (n_9));
NAND2_X1 slo__sro_c104 (.ZN (slo__sro_n183), .A1 (p_1[7]), .A2 (p_0[7]));
NOR2_X1 slo__sro_c105 (.ZN (slo__sro_n182), .A1 (p_1[7]), .A2 (p_0[7]));
OAI21_X1 slo__sro_c106 (.ZN (n_8), .A (slo__sro_n183), .B1 (slo__sro_n184), .B2 (slo__sro_n182));
XNOR2_X2 slo__sro_c107 (.ZN (slo__sro_n181), .A (p_1[7]), .B (p_0[7]));
XNOR2_X1 slo__sro_c108 (.ZN (p_2[7]), .A (slo__sro_n181), .B (n_7));
NAND2_X1 slo__sro_c118 (.ZN (slo__sro_n196), .A1 (p_1[4]), .A2 (p_0[4]));
NOR2_X1 slo__sro_c119 (.ZN (slo__sro_n195), .A1 (p_1[4]), .A2 (p_0[4]));
OAI21_X1 slo__sro_c120 (.ZN (n_5), .A (slo__sro_n196), .B1 (slo__sro_n197), .B2 (slo__sro_n195));
XNOR2_X1 slo__sro_c121 (.ZN (slo__sro_n194), .A (p_1[4]), .B (p_0[4]));
XNOR2_X1 slo__sro_c122 (.ZN (p_2[4]), .A (slo__sro_n194), .B (n_4));
NOR2_X1 slo__sro_c189 (.ZN (slo__sro_n293), .A1 (n_33), .A2 (p_0[30]));
NAND2_X1 slo__sro_c190 (.ZN (slo__sro_n292), .A1 (slo__sro_n293), .A2 (slo__sro_n294));
OR2_X1 slo__sro_c191 (.ZN (slo__sro_n291), .A1 (p_1[30]), .A2 (n_34));
OAI21_X1 slo__sro_c192 (.ZN (n_31), .A (slo__sro_n292), .B1 (n_32), .B2 (slo__sro_n291));
OAI21_X1 slo__sro_c201 (.ZN (slo__sro_n305), .A (n_21), .B1 (p_1[21]), .B2 (p_0[21]));
NAND2_X1 slo__sro_c202 (.ZN (slo__sro_n304), .A1 (slo__sro_n305), .A2 (slo__sro_n306));
XNOR2_X1 slo__sro_c203 (.ZN (slo__sro_n303), .A (n_21), .B (p_0[21]));
XNOR2_X1 slo__sro_c204 (.ZN (p_2[21]), .A (slo__sro_n303), .B (p_1[21]));
OAI21_X1 slo__sro_c213 (.ZN (slo__sro_n319), .A (n_20), .B1 (p_1[20]), .B2 (p_0[20]));
NAND2_X1 slo__sro_c214 (.ZN (n_21), .A1 (slo__sro_n319), .A2 (slo__sro_n320));
XNOR2_X1 slo__sro_c215 (.ZN (slo__sro_n318), .A (p_1[20]), .B (p_0[20]));
XNOR2_X1 slo__sro_c216 (.ZN (p_2[20]), .A (slo__sro_n318), .B (n_20));
AOI22_X1 slo__sro_c225 (.ZN (slo__sro_n332), .A1 (p_1[22]), .A2 (slo__sro_n304), .B1 (slo__sro_n304), .B2 (p_0[22]));
NAND2_X1 slo__sro_c226 (.ZN (n_23), .A1 (slo__sro_n332), .A2 (slo__sro_n333));
XNOR2_X1 slo__sro_c227 (.ZN (slo__sro_n331), .A (slo__sro_n304), .B (p_0[22]));
XNOR2_X1 slo__sro_c228 (.ZN (p_2[22]), .A (slo__sro_n331), .B (p_1[22]));
OAI21_X1 slo__sro_c237 (.ZN (slo__sro_n346), .A (n_25), .B1 (p_1[25]), .B2 (p_0[25]));
NAND2_X1 slo__sro_c238 (.ZN (slo__sro_n345), .A1 (slo__sro_n346), .A2 (slo__sro_n347));
XNOR2_X1 slo__sro_c239 (.ZN (slo__sro_n344), .A (p_1[25]), .B (p_0[25]));
XNOR2_X1 slo__sro_c240 (.ZN (p_2[25]), .A (slo__sro_n344), .B (n_25));
NAND2_X1 slo__sro_c299 (.ZN (slo__sro_n438), .A1 (p_1[23]), .A2 (p_0[23]));
NAND2_X1 slo__sro_c300 (.ZN (slo__sro_n437), .A1 (n_23), .A2 (p_0[23]));
NAND2_X1 slo__sro_c301 (.ZN (slo__sro_n436), .A1 (n_23), .A2 (p_1[23]));
NAND3_X1 slo__sro_c302 (.ZN (slo__sro_n435), .A1 (slo__sro_n436), .A2 (slo__sro_n438), .A3 (slo__sro_n437));
XNOR2_X2 slo__sro_c303 (.ZN (slo__sro_n434), .A (p_1[23]), .B (p_0[23]));
XNOR2_X1 slo__sro_c304 (.ZN (p_2[23]), .A (slo__sro_n434), .B (n_23));
XNOR2_X2 slo__mro_c317 (.ZN (p_2[1]), .A (p_1[1]), .B (slo__mro_n453));
NOR2_X1 slo__sro_c328 (.ZN (slo__sro_n471), .A1 (p_1[3]), .A2 (p_0[3]));
OAI21_X4 slo__sro_c329 (.ZN (n_4), .A (slo__sro_n472), .B1 (slo__sro_n473), .B2 (slo__sro_n471));
XNOR2_X1 slo__sro_c330 (.ZN (slo__sro_n470), .A (p_1[3]), .B (p_0[3]));
XNOR2_X1 slo__sro_c331 (.ZN (p_2[3]), .A (slo__sro_n470), .B (n_3));
NAND2_X1 slo__sro_c364 (.ZN (slo__sro_n512), .A1 (p_1[2]), .A2 (p_0[2]));
NOR2_X1 slo__sro_c365 (.ZN (slo__sro_n511), .A1 (p_1[2]), .A2 (p_0[2]));
NAND2_X1 slo__sro_c349 (.ZN (slo__sro_n494), .A1 (p_0[17]), .A2 (p_1[17]));
NAND2_X1 CLOCK_slo__sro_c696 (.ZN (CLOCK_slo__sro_n963), .A1 (p_1[24]), .A2 (p_0[24]));
NAND2_X1 slo__sro_c351 (.ZN (slo__sro_n492), .A1 (slo__sro_n493), .A2 (slo__sro_n494));
XNOR2_X1 slo__sro_c352 (.ZN (slo__sro_n491), .A (slo__sro_n114), .B (p_0[17]));
XNOR2_X1 slo__sro_c353 (.ZN (p_2[17]), .A (slo__sro_n491), .B (p_1[17]));
XNOR2_X1 slo__sro_c367 (.ZN (slo__sro_n510), .A (p_1[2]), .B (p_0[2]));
XNOR2_X1 slo__sro_c368 (.ZN (p_2[2]), .A (slo__sro_n131), .B (slo__sro_n510));
INV_X2 CLOCK_slo__sro_c530 (.ZN (CLOCK_slo__sro_n767), .A (p_1[0]));
NOR2_X2 CLOCK_slo__sro_c531 (.ZN (n_1), .A1 (CLOCK_slo__sro_n767), .A2 (CLOCK_slo__sro_n768));
XNOR2_X1 CLOCK_slo__sro_c532 (.ZN (p_2[0]), .A (p_1[0]), .B (CLOCK_slo__sro_n768));
NAND2_X1 CLOCK_slo__sro_c551 (.ZN (CLOCK_slo__sro_n789), .A1 (p_1[15]), .A2 (p_0[15]));
NOR2_X1 CLOCK_slo__sro_c552 (.ZN (CLOCK_slo__sro_n788), .A1 (p_1[15]), .A2 (p_0[15]));
OAI21_X1 CLOCK_slo__sro_c553 (.ZN (CLOCK_slo__sro_n787), .A (CLOCK_slo__sro_n789)
    , .B1 (CLOCK_slo__sro_n790), .B2 (CLOCK_slo__sro_n788));
XNOR2_X1 CLOCK_slo__sro_c554 (.ZN (CLOCK_slo__sro_n786), .A (p_1[15]), .B (p_0[15]));
XNOR2_X1 CLOCK_slo__sro_c555 (.ZN (p_2[15]), .A (n_15), .B (CLOCK_slo__sro_n786));
INV_X1 CLOCK_slo__sro_c634 (.ZN (CLOCK_slo__sro_n898), .A (p_0[31]));
XNOR2_X1 CLOCK_slo__sro_c635 (.ZN (p_2[31]), .A (n_31), .B (CLOCK_slo__sro_n898));
INV_X1 CLOCK_slo__sro_c653 (.ZN (CLOCK_slo__sro_n918), .A (p_0[17]));
NAND2_X1 CLOCK_slo__sro_c654 (.ZN (CLOCK_slo__sro_n917), .A1 (CLOCK_slo__sro_n919), .A2 (CLOCK_slo__sro_n918));
NAND2_X1 CLOCK_slo__sro_c655 (.ZN (slo__sro_n493), .A1 (slo__sro_n114), .A2 (CLOCK_slo__sro_n917));
NAND2_X1 CLOCK_slo__sro_c697 (.ZN (CLOCK_slo__sro_n962), .A1 (slo__sro_n435), .A2 (p_0[24]));
NAND2_X1 CLOCK_slo__sro_c698 (.ZN (CLOCK_slo__sro_n961), .A1 (p_1[24]), .A2 (slo__sro_n435));
NAND3_X1 CLOCK_slo__sro_c699 (.ZN (n_25), .A1 (CLOCK_slo__sro_n961), .A2 (CLOCK_slo__sro_n962), .A3 (CLOCK_slo__sro_n963));
XNOR2_X1 CLOCK_slo__sro_c700 (.ZN (CLOCK_slo__sro_n960), .A (p_1[24]), .B (p_0[24]));
XNOR2_X1 CLOCK_slo__sro_c701 (.ZN (p_2[24]), .A (CLOCK_slo__sro_n960), .B (slo__sro_n435));
INV_X1 CLOCK_slo__sro_c838 (.ZN (CLOCK_slo__sro_n1105), .A (n_12));
NAND2_X1 CLOCK_slo__sro_c839 (.ZN (CLOCK_slo__sro_n1104), .A1 (p_1[12]), .A2 (p_0[12]));
NOR2_X1 CLOCK_slo__sro_c840 (.ZN (CLOCK_slo__sro_n1103), .A1 (p_1[12]), .A2 (p_0[12]));
OAI21_X1 CLOCK_slo__sro_c841 (.ZN (CLOCK_slo__sro_n1102), .A (CLOCK_slo__sro_n1104)
    , .B1 (CLOCK_slo__sro_n1103), .B2 (CLOCK_slo__sro_n1105));
XNOR2_X1 CLOCK_slo__sro_c842 (.ZN (CLOCK_slo__sro_n1101), .A (p_1[12]), .B (p_0[12]));
XNOR2_X1 CLOCK_slo__sro_c843 (.ZN (p_2[12]), .A (CLOCK_slo__sro_n1101), .B (n_12));

endmodule //datapath__0_107

module datapath__0_106 (Multiplier, p_0, p_1);

output [31:0] p_1;
input [31:0] Multiplier;
input [31:0] p_0;
wire CLOCK_slo__sro_n1169;
wire slo__sro_n425;
wire CLOCK_slo__sro_n765;
wire n_1;
wire n_2;
wire n_4;
wire n_5;
wire n_6;
wire n_7;
wire n_10;
wire n_11;
wire n_12;
wire n_13;
wire n_14;
wire n_15;
wire CLOCK_slo__sro_n766;
wire n_17;
wire n_18;
wire n_19;
wire n_20;
wire n_22;
wire n_23;
wire n_25;
wire n_26;
wire slo__sro_n119;
wire n_28;
wire n_29;
wire n_32;
wire n_0;
wire n_34;
wire n_33;
wire n_31;
wire slo__sro_n106;
wire CLOCK_slo__sro_n1167;
wire slo__sro_n108;
wire slo__sro_n109;
wire slo__sro_n89;
wire slo__sro_n90;
wire slo__sro_n91;
wire slo__sro_n92;
wire slo__sro_n93;
wire slo__sro_n120;
wire slo__sro_n121;
wire slo__sro_n122;
wire slo__sro_n123;
wire slo__sro_n151;
wire slo__sro_n152;
wire slo__sro_n153;
wire slo__sro_n154;
wire slo__sro_n445;
wire slo__sro_n446;
wire CLOCK_slo__sro_n714;
wire slo__sro_n423;
wire slo__sro_n424;
wire slo__sro_n384;
wire slo__sro_n385;
wire slo__sro_n386;
wire slo__sro_n387;
wire slo__sro_n388;
wire slo__sro_n447;
wire slo__sro_n448;
wire slo__sro_n449;
wire slo__sro_n521;
wire slo__sro_n522;
wire slo__sro_n523;
wire slo__sro_n524;
wire slo__sro_n502;
wire slo__sro_n503;
wire slo__sro_n504;
wire slo__sro_n505;
wire slo__sro_n506;
wire CLOCK_opt_ipo_n654;
wire CLOCK_slo__mro_n696;
wire CLOCK_slo__sro_n715;
wire CLOCK_slo__sro_n716;
wire CLOCK_slo__sro_n717;
wire CLOCK_slo__sro_n1161;
wire CLOCK_slo__sro_n763;
wire CLOCK_slo__sro_n764;
wire CLOCK_slo__sro_n1168;
wire CLOCK_slo__sro_n804;
wire CLOCK_slo__sro_n805;
wire CLOCK_slo__sro_n806;
wire CLOCK_slo__sro_n850;
wire CLOCK_slo__sro_n851;
wire CLOCK_slo__sro_n852;
wire CLOCK_slo__sro_n853;
wire CLOCK_slo__sro_n854;
wire CLOCK_slo__sro_n935;
wire CLOCK_slo__sro_n936;
wire CLOCK_slo__sro_n937;
wire CLOCK_slo__sro_n938;
wire CLOCK_slo__sro_n939;


INV_X1 i_36 (.ZN (n_34), .A (Multiplier[30]));
INV_X1 i_35 (.ZN (n_33), .A (p_0[30]));
INV_X1 i_34 (.ZN (n_32), .A (CLOCK_slo__sro_n851));
OAI33_X1 i_33 (.ZN (n_31), .A1 (n_34), .A2 (p_0[30]), .A3 (n_32), .B1 (CLOCK_slo__sro_n851)
    , .B2 (n_33), .B3 (Multiplier[30]));
XOR2_X1 i_32 (.Z (p_1[31]), .A (Multiplier[31]), .B (n_31));
OAI22_X1 i_31 (.ZN (n_0), .A1 (n_34), .A2 (p_0[30]), .B1 (Multiplier[30]), .B2 (n_33));
XNOR2_X1 i_0 (.ZN (p_1[30]), .A (n_32), .B (n_0));
XNOR2_X1 CLOCK_slo__sro_c1006 (.ZN (CLOCK_slo__sro_n1167), .A (p_0[3]), .B (Multiplier[3]));
FA_X1 i_29 (.CO (n_29), .S (p_1[28]), .A (Multiplier[28]), .B (p_0[28]), .CI (n_28));
FA_X1 i_28 (.CO (n_28), .S (p_1[27]), .A (Multiplier[27]), .B (p_0[27]), .CI (slo__sro_n90));
NAND2_X1 slo__sro_c60 (.ZN (slo__sro_n122), .A1 (p_0[7]), .A2 (Multiplier[7]));
FA_X1 i_26 (.CO (n_26), .S (p_1[25]), .A (Multiplier[25]), .B (p_0[25]), .CI (n_25));
FA_X1 i_25 (.CO (n_25), .S (p_1[24]), .A (Multiplier[24]), .B (p_0[24]), .CI (slo__sro_n385));
INV_X1 CLOCK_slo__sro_c562 (.ZN (CLOCK_slo__sro_n717), .A (n_6));
FA_X1 i_23 (.CO (n_23), .S (p_1[22]), .A (Multiplier[22]), .B (p_0[22]), .CI (n_22));
FA_X1 i_22 (.CO (n_22), .S (p_1[21]), .A (Multiplier[21]), .B (p_0[21]), .CI (slo__sro_n446));
INV_X1 slo__sro_c417 (.ZN (slo__sro_n524), .A (n_14));
FA_X1 i_20 (.CO (n_20), .S (p_1[19]), .A (Multiplier[19]), .B (p_0[19]), .CI (n_19));
FA_X1 i_19 (.CO (n_19), .S (p_1[18]), .A (Multiplier[18]), .B (p_0[18]), .CI (n_18));
FA_X1 i_18 (.CO (n_18), .S (p_1[17]), .A (Multiplier[17]), .B (p_0[17]), .CI (n_17));
FA_X1 i_17 (.CO (n_17), .S (p_1[16]), .A (Multiplier[16]), .B (p_0[16]), .CI (slo__sro_n503));
XNOR2_X1 CLOCK_slo__sro_c619 (.ZN (p_1[9]), .A (CLOCK_slo__sro_n763), .B (CLOCK_slo__sro_n936));
XNOR2_X1 CLOCK_slo__sro_c618 (.ZN (CLOCK_slo__sro_n763), .A (p_0[9]), .B (Multiplier[9]));
NOR2_X1 slo__sro_c348 (.ZN (slo__sro_n447), .A1 (p_0[20]), .A2 (Multiplier[20]));
FA_X1 i_13 (.CO (n_13), .S (p_1[12]), .A (Multiplier[12]), .B (p_0[12]), .CI (n_12));
FA_X1 i_12 (.CO (n_12), .S (p_1[11]), .A (Multiplier[11]), .B (p_0[11]), .CI (n_11));
FA_X1 i_11 (.CO (n_11), .S (p_1[10]), .A (Multiplier[10]), .B (p_0[10]), .CI (n_10));
NOR2_X2 CLOCK_slo__sro_c999 (.ZN (CLOCK_slo__sro_n1161), .A1 (p_0[1]), .A2 (Multiplier[1]));
INV_X1 slo__sro_c86 (.ZN (slo__sro_n154), .A (n_13));
NAND2_X1 CLOCK_slo__sro_c1003 (.ZN (CLOCK_slo__sro_n1169), .A1 (slo__sro_n423), .A2 (Multiplier[3]));
FA_X1 i_6 (.CO (n_6), .S (p_1[5]), .A (Multiplier[5]), .B (p_0[5]), .CI (n_5));
FA_X1 i_5 (.CO (n_5), .S (p_1[4]), .A (Multiplier[4]), .B (p_0[4]), .CI (n_4));
INV_X1 slo__sro_c346 (.ZN (slo__sro_n449), .A (n_20));
INV_X1 slo__sro_c59 (.ZN (slo__sro_n123), .A (n_7));
HA_X1 i_1 (.CO (n_1), .S (p_1[0]), .A (Multiplier[0]), .B (p_0[0]));
INV_X1 slo__sro_c45 (.ZN (slo__sro_n109), .A (n_1));
NAND2_X1 slo__sro_c46 (.ZN (slo__sro_n108), .A1 (p_0[1]), .A2 (Multiplier[1]));
NAND2_X1 CLOCK_slo__sro_c1005 (.ZN (n_4), .A1 (CLOCK_slo__sro_n1168), .A2 (CLOCK_slo__sro_n1169));
OAI21_X2 slo__sro_c48 (.ZN (n_2), .A (slo__sro_n108), .B1 (CLOCK_slo__sro_n1161), .B2 (slo__sro_n109));
XNOR2_X2 slo__sro_c49 (.ZN (slo__sro_n106), .A (p_0[1]), .B (Multiplier[1]));
XNOR2_X2 slo__sro_c50 (.ZN (p_1[1]), .A (slo__sro_n106), .B (n_1));
INV_X1 slo__sro_c31 (.ZN (slo__sro_n93), .A (n_26));
NAND2_X1 slo__sro_c32 (.ZN (slo__sro_n92), .A1 (p_0[26]), .A2 (Multiplier[26]));
NOR2_X1 slo__sro_c33 (.ZN (slo__sro_n91), .A1 (p_0[26]), .A2 (Multiplier[26]));
OAI21_X1 slo__sro_c34 (.ZN (slo__sro_n90), .A (slo__sro_n92), .B1 (slo__sro_n93), .B2 (slo__sro_n91));
XNOR2_X1 slo__sro_c35 (.ZN (slo__sro_n89), .A (p_0[26]), .B (Multiplier[26]));
XNOR2_X1 slo__sro_c36 (.ZN (p_1[26]), .A (slo__sro_n89), .B (n_26));
NOR2_X1 slo__sro_c61 (.ZN (slo__sro_n121), .A1 (p_0[7]), .A2 (Multiplier[7]));
OAI21_X1 slo__sro_c62 (.ZN (slo__sro_n120), .A (slo__sro_n122), .B1 (slo__sro_n123), .B2 (slo__sro_n121));
XNOR2_X1 slo__sro_c63 (.ZN (slo__sro_n119), .A (p_0[7]), .B (Multiplier[7]));
XNOR2_X1 slo__sro_c64 (.ZN (p_1[7]), .A (n_7), .B (slo__sro_n119));
NAND2_X1 slo__sro_c87 (.ZN (slo__sro_n153), .A1 (p_0[13]), .A2 (Multiplier[13]));
NOR2_X1 slo__sro_c88 (.ZN (slo__sro_n152), .A1 (p_0[13]), .A2 (Multiplier[13]));
OAI21_X2 slo__sro_c89 (.ZN (n_14), .A (slo__sro_n153), .B1 (slo__sro_n154), .B2 (slo__sro_n152));
XNOR2_X1 slo__sro_c90 (.ZN (slo__sro_n151), .A (p_0[13]), .B (Multiplier[13]));
XNOR2_X1 slo__sro_c91 (.ZN (p_1[13]), .A (n_13), .B (slo__sro_n151));
OAI21_X1 slo__sro_c349 (.ZN (slo__sro_n446), .A (slo__sro_n448), .B1 (slo__sro_n449), .B2 (slo__sro_n447));
NAND2_X1 slo__sro_c330 (.ZN (slo__sro_n425), .A1 (CLOCK_opt_ipo_n654), .A2 (Multiplier[2]));
INV_X1 CLOCK_slo__sro_c681 (.ZN (CLOCK_slo__sro_n854), .A (n_29));
NAND2_X2 slo__sro_c332 (.ZN (slo__sro_n423), .A1 (slo__sro_n424), .A2 (slo__sro_n425));
AOI22_X2 CLOCK_slo__sro_c1004 (.ZN (CLOCK_slo__sro_n1168), .A1 (slo__sro_n423), .A2 (p_0[3])
    , .B1 (p_0[3]), .B2 (Multiplier[3]));
INV_X1 slo__sro_c293 (.ZN (slo__sro_n388), .A (n_23));
NAND2_X1 slo__sro_c294 (.ZN (slo__sro_n387), .A1 (p_0[23]), .A2 (Multiplier[23]));
NOR2_X1 slo__sro_c295 (.ZN (slo__sro_n386), .A1 (p_0[23]), .A2 (Multiplier[23]));
OAI21_X1 slo__sro_c296 (.ZN (slo__sro_n385), .A (slo__sro_n387), .B1 (slo__sro_n388), .B2 (slo__sro_n386));
XNOR2_X1 slo__sro_c297 (.ZN (slo__sro_n384), .A (p_0[23]), .B (Multiplier[23]));
XNOR2_X1 slo__sro_c298 (.ZN (p_1[23]), .A (slo__sro_n384), .B (n_23));
NAND2_X1 slo__sro_c347 (.ZN (slo__sro_n448), .A1 (p_0[20]), .A2 (Multiplier[20]));
XNOR2_X2 slo__sro_c350 (.ZN (slo__sro_n445), .A (p_0[20]), .B (Multiplier[20]));
XNOR2_X2 slo__sro_c351 (.ZN (p_1[20]), .A (n_20), .B (slo__sro_n445));
NAND2_X1 slo__sro_c418 (.ZN (slo__sro_n523), .A1 (p_0[14]), .A2 (Multiplier[14]));
NOR2_X1 slo__sro_c419 (.ZN (slo__sro_n522), .A1 (p_0[14]), .A2 (Multiplier[14]));
OAI21_X2 slo__sro_c420 (.ZN (n_15), .A (slo__sro_n523), .B1 (slo__sro_n524), .B2 (slo__sro_n522));
XNOR2_X1 slo__sro_c421 (.ZN (slo__sro_n521), .A (p_0[14]), .B (Multiplier[14]));
XNOR2_X1 slo__sro_c422 (.ZN (p_1[14]), .A (slo__sro_n521), .B (n_14));
INV_X2 slo__sro_c401 (.ZN (slo__sro_n506), .A (n_15));
NAND2_X1 slo__sro_c402 (.ZN (slo__sro_n505), .A1 (p_0[15]), .A2 (Multiplier[15]));
NOR2_X1 slo__sro_c403 (.ZN (slo__sro_n504), .A1 (p_0[15]), .A2 (Multiplier[15]));
OAI21_X1 slo__sro_c404 (.ZN (slo__sro_n503), .A (slo__sro_n505), .B1 (slo__sro_n506), .B2 (slo__sro_n504));
XNOR2_X1 slo__sro_c405 (.ZN (slo__sro_n502), .A (p_0[15]), .B (Multiplier[15]));
XNOR2_X1 slo__sro_c406 (.ZN (p_1[15]), .A (slo__sro_n502), .B (n_15));
INV_X4 CLOCK_opt_ipo_c528 (.ZN (CLOCK_opt_ipo_n654), .A (p_0[2]));
XNOR2_X2 CLOCK_slo__mro_c541 (.ZN (CLOCK_slo__mro_n696), .A (CLOCK_opt_ipo_n654), .B (Multiplier[2]));
XNOR2_X2 CLOCK_slo__mro_c542 (.ZN (p_1[2]), .A (CLOCK_slo__mro_n696), .B (n_2));
NAND2_X1 CLOCK_slo__sro_c563 (.ZN (CLOCK_slo__sro_n716), .A1 (p_0[6]), .A2 (Multiplier[6]));
NOR2_X1 CLOCK_slo__sro_c564 (.ZN (CLOCK_slo__sro_n715), .A1 (p_0[6]), .A2 (Multiplier[6]));
OAI21_X1 CLOCK_slo__sro_c565 (.ZN (n_7), .A (CLOCK_slo__sro_n716), .B1 (CLOCK_slo__sro_n717), .B2 (CLOCK_slo__sro_n715));
XNOR2_X2 CLOCK_slo__sro_c566 (.ZN (CLOCK_slo__sro_n714), .A (p_0[6]), .B (Multiplier[6]));
XNOR2_X1 CLOCK_slo__sro_c567 (.ZN (p_1[6]), .A (CLOCK_slo__sro_n714), .B (n_6));
INV_X2 CLOCK_slo__sro_c614 (.ZN (CLOCK_slo__sro_n766), .A (CLOCK_slo__sro_n936));
NAND2_X1 CLOCK_slo__sro_c615 (.ZN (CLOCK_slo__sro_n765), .A1 (p_0[9]), .A2 (Multiplier[9]));
NOR2_X1 CLOCK_slo__sro_c616 (.ZN (CLOCK_slo__sro_n764), .A1 (p_0[9]), .A2 (Multiplier[9]));
OAI21_X2 CLOCK_slo__sro_c617 (.ZN (n_10), .A (CLOCK_slo__sro_n765), .B1 (CLOCK_slo__sro_n766), .B2 (CLOCK_slo__sro_n764));
INV_X1 CLOCK_slo__sro_c644 (.ZN (CLOCK_slo__sro_n806), .A (CLOCK_opt_ipo_n654));
INV_X1 CLOCK_slo__sro_c645 (.ZN (CLOCK_slo__sro_n805), .A (Multiplier[2]));
NAND2_X1 CLOCK_slo__sro_c646 (.ZN (CLOCK_slo__sro_n804), .A1 (CLOCK_slo__sro_n806), .A2 (CLOCK_slo__sro_n805));
NAND2_X2 CLOCK_slo__sro_c647 (.ZN (slo__sro_n424), .A1 (n_2), .A2 (CLOCK_slo__sro_n804));
NAND2_X1 CLOCK_slo__sro_c682 (.ZN (CLOCK_slo__sro_n853), .A1 (p_0[29]), .A2 (Multiplier[29]));
NOR2_X1 CLOCK_slo__sro_c683 (.ZN (CLOCK_slo__sro_n852), .A1 (p_0[29]), .A2 (Multiplier[29]));
OAI21_X1 CLOCK_slo__sro_c684 (.ZN (CLOCK_slo__sro_n851), .A (CLOCK_slo__sro_n853)
    , .B1 (CLOCK_slo__sro_n854), .B2 (CLOCK_slo__sro_n852));
XNOR2_X1 CLOCK_slo__sro_c685 (.ZN (CLOCK_slo__sro_n850), .A (p_0[29]), .B (Multiplier[29]));
XNOR2_X1 CLOCK_slo__sro_c686 (.ZN (p_1[29]), .A (CLOCK_slo__sro_n850), .B (n_29));
XNOR2_X1 CLOCK_slo__sro_c1007 (.ZN (p_1[3]), .A (CLOCK_slo__sro_n1167), .B (slo__sro_n423));
NAND2_X1 CLOCK_slo__sro_c748 (.ZN (CLOCK_slo__sro_n939), .A1 (p_0[8]), .A2 (Multiplier[8]));
NAND2_X1 CLOCK_slo__sro_c749 (.ZN (CLOCK_slo__sro_n938), .A1 (slo__sro_n120), .A2 (Multiplier[8]));
NAND2_X1 CLOCK_slo__sro_c750 (.ZN (CLOCK_slo__sro_n937), .A1 (slo__sro_n120), .A2 (p_0[8]));
NAND3_X2 CLOCK_slo__sro_c751 (.ZN (CLOCK_slo__sro_n936), .A1 (CLOCK_slo__sro_n938)
    , .A2 (CLOCK_slo__sro_n937), .A3 (CLOCK_slo__sro_n939));
XNOR2_X2 CLOCK_slo__sro_c752 (.ZN (CLOCK_slo__sro_n935), .A (p_0[8]), .B (Multiplier[8]));
XNOR2_X1 CLOCK_slo__sro_c753 (.ZN (p_1[8]), .A (CLOCK_slo__sro_n935), .B (slo__sro_n120));

endmodule //datapath__0_106

module datapath__0_102 (p_0_9_PP_0, opt_ipoPP_2, p_0, p_1, p_2);

output [31:0] p_2;
input [31:0] p_0;
input [31:0] p_1;
input p_0_9_PP_0;
input opt_ipoPP_2;
wire n_6;
wire n_7;
wire n_8;
wire n_10;
wire n_12;
wire n_14;
wire CLOCK_slo__sro_n932;
wire n_16;
wire n_17;
wire n_18;
wire n_19;
wire n_20;
wire n_21;
wire n_22;
wire n_23;
wire n_24;
wire n_25;
wire n_26;
wire n_27;
wire n_28;
wire n_29;
wire n_30;
wire n_32;
wire n_0;
wire n_34;
wire n_33;
wire slo__sro_n65;
wire slo__sro_n66;
wire slo__sro_n68;
wire CLOCK_slo__sro_n931;
wire slo__sro_n81;
wire slo__sro_n82;
wire slo__sro_n83;
wire slo__sro_n84;
wire slo__sro_n99;
wire slo__sro_n100;
wire slo__sro_n101;
wire slo__sro_n102;
wire slo__sro_n103;
wire slo__sro_n131;
wire slo__sro_n132;
wire slo__sro_n133;
wire slo__sro_n134;
wire slo__sro_n135;
wire slo__sro_n150;
wire slo__sro_n151;
wire slo__sro_n152;
wire slo__sro_n153;
wire slo__sro_n167;
wire slo__sro_n168;
wire slo__sro_n169;
wire slo__sro_n170;
wire slo__sro_n171;
wire slo__sro_n187;
wire slo__sro_n188;
wire slo__sro_n189;
wire slo__sro_n190;
wire slo__sro_n191;
wire slo__sro_n208;
wire slo__sro_n209;
wire slo__sro_n210;
wire slo__sro_n211;
wire slo__sro_n212;
wire slo__sro_n375;
wire slo__sro_n376;
wire slo__sro_n377;
wire slo__sro_n427;
wire slo__sro_n428;
wire slo__sro_n429;
wire slo__sro_n430;
wire CLOCK_slo__mro_n891;
wire CLOCK_slo__sro_n933;
wire CLOCK_slo__sro_n934;
wire CLOCK_slo__sro_n945;
wire CLOCK_slo__sro_n946;
wire CLOCK_slo__sro_n947;
wire CLOCK_slo__sro_n948;
wire CLOCK_slo__sro_n949;
wire CLOCK_slo__sro_n950;
wire CLOCK_slo__sro_n1043;
wire CLOCK_slo__sro_n1044;
wire CLOCK_slo__sro_n1045;
wire CLOCK_slo__sro_n1046;
wire CLOCK_slo__sro_n1047;
wire CLOCK_slo__sro_n990;
wire CLOCK_slo__sro_n991;
wire CLOCK_slo__sro_n992;
wire CLOCK_slo__sro_n993;
wire CLOCK_slo__sro_n1145;
wire CLOCK_slo__sro_n1146;
wire CLOCK_slo__sro_n1147;
wire CLOCK_slo__sro_n1148;


INV_X1 i_36 (.ZN (n_34), .A (p_0[30]));
INV_X1 i_35 (.ZN (n_33), .A (p_1[30]));
INV_X1 i_34 (.ZN (n_32), .A (n_30));
INV_X2 CLOCK_slo__sro_c763 (.ZN (CLOCK_slo__sro_n1148), .A (n_18));
XOR2_X1 i_32 (.Z (p_2[31]), .A (p_0[31]), .B (CLOCK_slo__sro_n1043));
OAI22_X1 i_31 (.ZN (n_0), .A1 (n_34), .A2 (p_1[30]), .B1 (p_0[30]), .B2 (n_33));
XNOR2_X1 i_0 (.ZN (p_2[30]), .A (n_32), .B (n_0));
FA_X1 i_30 (.CO (n_30), .S (p_2[29]), .A (p_0[29]), .B (p_1[29]), .CI (n_29));
FA_X1 i_29 (.CO (n_29), .S (p_2[28]), .A (p_0[28]), .B (p_1[28]), .CI (n_28));
FA_X1 i_28 (.CO (n_28), .S (p_2[27]), .A (p_0[27]), .B (p_1[27]), .CI (n_27));
FA_X1 i_27 (.CO (n_27), .S (p_2[26]), .A (p_0[26]), .B (p_1[26]), .CI (n_26));
FA_X1 i_26 (.CO (n_26), .S (p_2[25]), .A (p_0[25]), .B (p_1[25]), .CI (n_25));
FA_X1 i_25 (.CO (n_25), .S (p_2[24]), .A (p_0[24]), .B (p_1[24]), .CI (n_24));
FA_X1 i_24 (.CO (n_24), .S (p_2[23]), .A (p_0[23]), .B (p_1[23]), .CI (n_23));
FA_X1 i_23 (.CO (n_23), .S (p_2[22]), .A (p_0[22]), .B (p_1[22]), .CI (n_22));
FA_X1 i_22 (.CO (n_22), .S (p_2[21]), .A (p_0[21]), .B (p_1[21]), .CI (n_21));
NOR2_X1 CLOCK_slo__sro_c765 (.ZN (CLOCK_slo__sro_n1146), .A1 (p_1[18]), .A2 (p_0[18]));
FA_X1 i_20 (.CO (n_20), .S (p_2[19]), .A (p_0[19]), .B (p_1[19]), .CI (n_19));
FA_X1 i_18 (.CO (n_18), .S (p_2[17]), .A (p_0[17]), .B (p_1[17]), .CI (n_17));
FA_X1 i_17 (.CO (n_17), .S (p_2[16]), .A (p_0[16]), .B (p_1[16]), .CI (n_16));
FA_X1 i_16 (.CO (n_16), .S (p_2[15]), .A (p_0[15]), .B (p_1[15]), .CI (slo__sro_n66));
INV_X2 slo__sro_c15 (.ZN (slo__sro_n84), .A (slo__sro_n209));
FA_X1 i_14 (.CO (n_14), .S (p_2[13]), .A (p_0[13]), .B (p_1[13]), .CI (slo__sro_n100));
INV_X2 slo__sro_c58 (.ZN (slo__sro_n135), .A (n_10));
INV_X1 CLOCK_slo__sro_c652 (.ZN (CLOCK_slo__sro_n1047), .A (n_30));
INV_X1 slo__sro_c74 (.ZN (slo__sro_n153), .A (slo__sro_n168));
INV_X1 slo__sro_c90 (.ZN (slo__sro_n171), .A (n_8));
INV_X2 slo__sro_c107 (.ZN (slo__sro_n191), .A (slo__sro_n81));
FA_X1 i_8 (.CO (n_8), .S (p_2[7]), .A (p_0[7]), .B (p_1[7]), .CI (n_7));
FA_X1 i_7 (.CO (n_7), .S (p_2[6]), .A (p_0[6]), .B (p_1[6]), .CI (n_6));
FA_X1 i_6 (.CO (n_6), .S (p_2[5]), .A (p_0[5]), .B (p_1[5]), .CI (slo__sro_n428));
XNOR2_X2 CLOCK_slo__mro_c481 (.ZN (p_2[2]), .A (CLOCK_slo__mro_n891), .B (slo__sro_n209));
NAND2_X2 slo__sro_c126 (.ZN (slo__sro_n212), .A1 (p_1[1]), .A2 (p_0[1]));
INV_X1 slo__sro_c31 (.ZN (slo__sro_n103), .A (n_12));
INV_X1 slo__sro_c245 (.ZN (slo__sro_n377), .A (p_0[0]));
NAND2_X1 slo__sro_c295 (.ZN (slo__sro_n430), .A1 (slo__sro_n188), .A2 (p_0[4]));
NAND2_X1 slo__sro_c3 (.ZN (slo__sro_n68), .A1 (p_1[14]), .A2 (p_0[14]));
INV_X1 CLOCK_slo__sro_c544 (.ZN (CLOCK_slo__sro_n950), .A (p_0[11]));
NAND2_X1 slo__sro_c5 (.ZN (slo__sro_n66), .A1 (CLOCK_slo__sro_n931), .A2 (slo__sro_n68));
XNOR2_X1 slo__sro_c6 (.ZN (slo__sro_n65), .A (p_1[14]), .B (p_0[14]));
XNOR2_X1 slo__sro_c7 (.ZN (p_2[14]), .A (slo__sro_n65), .B (n_14));
NAND2_X1 slo__sro_c16 (.ZN (slo__sro_n83), .A1 (p_1[2]), .A2 (p_0[2]));
NOR2_X2 slo__sro_c17 (.ZN (slo__sro_n82), .A1 (p_1[2]), .A2 (p_0[2]));
OAI21_X4 slo__sro_c18 (.ZN (slo__sro_n81), .A (slo__sro_n83), .B1 (slo__sro_n82), .B2 (slo__sro_n84));
INV_X1 CLOCK_slo__sro_c532 (.ZN (CLOCK_slo__sro_n934), .A (p_1[14]));
INV_X1 CLOCK_slo__sro_c533 (.ZN (CLOCK_slo__sro_n933), .A (p_0[14]));
NAND2_X1 slo__sro_c32 (.ZN (slo__sro_n102), .A1 (p_1[12]), .A2 (p_0[12]));
NOR2_X1 slo__sro_c33 (.ZN (slo__sro_n101), .A1 (p_1[12]), .A2 (p_0[12]));
OAI21_X1 slo__sro_c34 (.ZN (slo__sro_n100), .A (slo__sro_n102), .B1 (slo__sro_n103), .B2 (slo__sro_n101));
XNOR2_X1 slo__sro_c35 (.ZN (slo__sro_n99), .A (p_1[12]), .B (p_0[12]));
XNOR2_X1 slo__sro_c36 (.ZN (p_2[12]), .A (n_12), .B (slo__sro_n99));
NAND2_X1 slo__sro_c59 (.ZN (slo__sro_n134), .A1 (p_1[10]), .A2 (p_0[10]));
NOR2_X1 slo__sro_c60 (.ZN (slo__sro_n133), .A1 (p_1[10]), .A2 (p_0[10]));
OAI21_X2 slo__sro_c61 (.ZN (slo__sro_n132), .A (slo__sro_n134), .B1 (slo__sro_n135), .B2 (slo__sro_n133));
XNOR2_X1 slo__sro_c62 (.ZN (slo__sro_n131), .A (p_1[10]), .B (p_0[10]));
XNOR2_X1 slo__sro_c63 (.ZN (p_2[10]), .A (n_10), .B (slo__sro_n131));
NAND2_X1 slo__sro_c75 (.ZN (slo__sro_n152), .A1 (p_1[9]), .A2 (p_0[9]));
NOR2_X1 slo__sro_c76 (.ZN (slo__sro_n151), .A1 (p_1[9]), .A2 (p_0[9]));
OAI21_X2 slo__sro_c77 (.ZN (n_10), .A (slo__sro_n152), .B1 (slo__sro_n153), .B2 (slo__sro_n151));
XNOR2_X1 slo__sro_c78 (.ZN (slo__sro_n150), .A (p_1[9]), .B (p_0_9_PP_0));
XNOR2_X2 slo__sro_c79 (.ZN (p_2[9]), .A (slo__sro_n168), .B (slo__sro_n150));
NAND2_X1 slo__sro_c91 (.ZN (slo__sro_n170), .A1 (p_1[8]), .A2 (p_0[8]));
NOR2_X1 slo__sro_c92 (.ZN (slo__sro_n169), .A1 (p_1[8]), .A2 (p_0[8]));
OAI21_X2 slo__sro_c93 (.ZN (slo__sro_n168), .A (slo__sro_n170), .B1 (slo__sro_n171), .B2 (slo__sro_n169));
XNOR2_X1 slo__sro_c94 (.ZN (slo__sro_n167), .A (p_1[8]), .B (p_0[8]));
XNOR2_X1 slo__sro_c95 (.ZN (p_2[8]), .A (slo__sro_n167), .B (n_8));
NAND2_X1 slo__sro_c108 (.ZN (slo__sro_n190), .A1 (p_1[3]), .A2 (p_0[3]));
NOR2_X4 slo__sro_c109 (.ZN (slo__sro_n189), .A1 (p_1[3]), .A2 (p_0[3]));
OAI21_X4 slo__sro_c110 (.ZN (slo__sro_n188), .A (slo__sro_n190), .B1 (slo__sro_n191), .B2 (slo__sro_n189));
XNOR2_X2 slo__sro_c111 (.ZN (slo__sro_n187), .A (p_1[3]), .B (p_0[3]));
XNOR2_X2 slo__sro_c112 (.ZN (p_2[3]), .A (slo__sro_n187), .B (slo__sro_n81));
NAND2_X1 slo__sro_c127 (.ZN (slo__sro_n211), .A1 (slo__sro_n375), .A2 (p_0[1]));
NAND2_X2 slo__sro_c128 (.ZN (slo__sro_n210), .A1 (slo__sro_n375), .A2 (p_1[1]));
NAND3_X4 slo__sro_c129 (.ZN (slo__sro_n209), .A1 (slo__sro_n210), .A2 (slo__sro_n212), .A3 (slo__sro_n211));
XNOR2_X1 slo__sro_c130 (.ZN (slo__sro_n208), .A (slo__sro_n375), .B (p_0[1]));
XNOR2_X1 slo__sro_c131 (.ZN (p_2[1]), .A (slo__sro_n208), .B (p_1[1]));
NAND2_X2 slo__sro_c246 (.ZN (slo__sro_n376), .A1 (p_1[0]), .A2 (p_0[0]));
INV_X2 slo__sro_c247 (.ZN (slo__sro_n375), .A (slo__sro_n376));
XNOR2_X1 slo__sro_c248 (.ZN (p_2[0]), .A (opt_ipoPP_2), .B (slo__sro_n377));
AOI22_X1 slo__sro_c296 (.ZN (slo__sro_n429), .A1 (slo__sro_n188), .A2 (p_1[4]), .B1 (p_1[4]), .B2 (p_0[4]));
NAND2_X1 slo__sro_c297 (.ZN (slo__sro_n428), .A1 (slo__sro_n429), .A2 (slo__sro_n430));
XNOR2_X1 slo__sro_c298 (.ZN (slo__sro_n427), .A (p_1[4]), .B (p_0[4]));
XNOR2_X1 slo__sro_c299 (.ZN (p_2[4]), .A (slo__sro_n427), .B (slo__sro_n188));
NAND2_X1 CLOCK_slo__sro_c534 (.ZN (CLOCK_slo__sro_n932), .A1 (CLOCK_slo__sro_n933), .A2 (CLOCK_slo__sro_n934));
XNOR2_X2 CLOCK_slo__mro_c480 (.ZN (CLOCK_slo__mro_n891), .A (p_1[2]), .B (p_0[2]));
NAND2_X1 CLOCK_slo__sro_c535 (.ZN (CLOCK_slo__sro_n931), .A1 (n_14), .A2 (CLOCK_slo__sro_n932));
INV_X1 CLOCK_slo__sro_c545 (.ZN (CLOCK_slo__sro_n949), .A (p_1[11]));
NAND2_X1 CLOCK_slo__sro_c546 (.ZN (CLOCK_slo__sro_n948), .A1 (p_1[11]), .A2 (p_0[11]));
NAND2_X1 CLOCK_slo__sro_c547 (.ZN (CLOCK_slo__sro_n947), .A1 (CLOCK_slo__sro_n949), .A2 (CLOCK_slo__sro_n950));
NAND2_X2 CLOCK_slo__sro_c548 (.ZN (CLOCK_slo__sro_n946), .A1 (slo__sro_n132), .A2 (CLOCK_slo__sro_n947));
NAND2_X1 CLOCK_slo__sro_c549 (.ZN (n_12), .A1 (CLOCK_slo__sro_n946), .A2 (CLOCK_slo__sro_n948));
XNOR2_X1 CLOCK_slo__sro_c550 (.ZN (CLOCK_slo__sro_n945), .A (p_1[11]), .B (p_0[11]));
XNOR2_X1 CLOCK_slo__sro_c551 (.ZN (p_2[11]), .A (slo__sro_n132), .B (CLOCK_slo__sro_n945));
NOR2_X1 CLOCK_slo__sro_c653 (.ZN (CLOCK_slo__sro_n1046), .A1 (n_33), .A2 (p_0[30]));
NAND2_X1 CLOCK_slo__sro_c654 (.ZN (CLOCK_slo__sro_n1045), .A1 (CLOCK_slo__sro_n1046), .A2 (CLOCK_slo__sro_n1047));
OR2_X1 CLOCK_slo__sro_c655 (.ZN (CLOCK_slo__sro_n1044), .A1 (p_1[30]), .A2 (n_34));
OAI21_X1 CLOCK_slo__sro_c656 (.ZN (CLOCK_slo__sro_n1043), .A (CLOCK_slo__sro_n1045)
    , .B1 (n_32), .B2 (CLOCK_slo__sro_n1044));
NAND2_X1 CLOCK_slo__sro_c764 (.ZN (CLOCK_slo__sro_n1147), .A1 (p_1[18]), .A2 (p_0[18]));
INV_X2 CLOCK_slo__sro_c592 (.ZN (CLOCK_slo__sro_n993), .A (n_20));
NAND2_X1 CLOCK_slo__sro_c593 (.ZN (CLOCK_slo__sro_n992), .A1 (p_1[20]), .A2 (p_0[20]));
NOR2_X2 CLOCK_slo__sro_c594 (.ZN (CLOCK_slo__sro_n991), .A1 (p_1[20]), .A2 (p_0[20]));
OAI21_X2 CLOCK_slo__sro_c595 (.ZN (n_21), .A (CLOCK_slo__sro_n992), .B1 (CLOCK_slo__sro_n991), .B2 (CLOCK_slo__sro_n993));
XNOR2_X1 CLOCK_slo__sro_c596 (.ZN (CLOCK_slo__sro_n990), .A (p_1[20]), .B (p_0[20]));
XNOR2_X1 CLOCK_slo__sro_c597 (.ZN (p_2[20]), .A (CLOCK_slo__sro_n990), .B (n_20));
OAI21_X2 CLOCK_slo__sro_c766 (.ZN (n_19), .A (CLOCK_slo__sro_n1147), .B1 (CLOCK_slo__sro_n1146), .B2 (CLOCK_slo__sro_n1148));
XNOR2_X1 CLOCK_slo__sro_c767 (.ZN (CLOCK_slo__sro_n1145), .A (p_1[18]), .B (p_0[18]));
XNOR2_X1 CLOCK_slo__sro_c768 (.ZN (p_2[18]), .A (CLOCK_slo__sro_n1145), .B (n_18));

endmodule //datapath__0_102

module datapath__0_101 (opt_ipoPP_3, Multiplier, p_0, p_1);

output [31:0] p_1;
input [31:0] Multiplier;
input [31:0] p_0;
input opt_ipoPP_3;
wire n_1;
wire n_3;
wire n_4;
wire n_6;
wire slo__sro_n745;
wire n_8;
wire n_9;
wire n_10;
wire CLOCK_slo__sro_n1405;
wire n_12;
wire n_13;
wire n_15;
wire CLOCK_slo__sro_n1221;
wire n_18;
wire n_19;
wire n_21;
wire n_22;
wire n_23;
wire n_24;
wire n_25;
wire n_26;
wire n_27;
wire n_28;
wire n_29;
wire n_30;
wire n_32;
wire n_0;
wire n_34;
wire n_33;
wire n_31;
wire slo__sro_n63;
wire slo__sro_n64;
wire slo__sro_n65;
wire slo__sro_n66;
wire slo__sro_n78;
wire slo__sro_n79;
wire slo__sro_n80;
wire slo__sro_n81;
wire slo__sro_n82;
wire slo__sro_n96;
wire slo__sro_n97;
wire slo__sro_n98;
wire slo__sro_n99;
wire slo__sro_n114;
wire slo__sro_n115;
wire slo__sro_n116;
wire slo__sro_n117;
wire slo__sro_n127;
wire slo__sro_n128;
wire slo__sro_n129;
wire slo__n168;
wire slo__sro_n147;
wire slo__sro_n148;
wire slo__sro_n214;
wire slo__sro_n215;
wire slo__sro_n216;
wire slo__sro_n217;
wire slo__sro_n855;
wire slo__sro_n746;
wire slo__sro_n747;
wire slo__sro_n748;
wire slo__sro_n760;
wire slo__sro_n761;
wire slo__sro_n762;
wire slo__sro_n763;
wire slo__sro_n777;
wire slo__sro_n778;
wire slo__sro_n779;
wire slo__sro_n780;
wire slo__sro_n781;
wire slo__sro_n827;
wire slo__sro_n828;
wire slo__sro_n829;
wire slo__sro_n830;
wire slo__sro_n831;
wire slo__mro_n844;
wire slo__sro_n856;
wire slo__sro_n857;
wire CLOCK_slo__sro_n1185;
wire CLOCK_slo__sro_n1186;
wire CLOCK_slo__sro_n1187;
wire CLOCK_slo__sro_n1218;
wire CLOCK_slo__sro_n1219;
wire CLOCK_slo__sro_n1220;
wire CLOCK_slo__sro_n1208;
wire CLOCK_slo__sro_n1209;
wire CLOCK_slo__sro_n1210;
wire slo__sro_n918;
wire slo__sro_n919;
wire slo__sro_n920;
wire slo__sro_n921;
wire slo__sro_n922;
wire CLOCK_slo__sro_n1222;
wire CLOCK_slo__sro_n1401;
wire CLOCK_slo__sro_n1255;
wire CLOCK_slo__sro_n1256;
wire CLOCK_slo__sro_n1257;
wire CLOCK_slo__sro_n1258;
wire CLOCK_slo__sro_n1402;
wire CLOCK_slo__sro_n1403;
wire CLOCK_slo__sro_n1404;
wire CLOCK_slo__sro_n1315;
wire CLOCK_slo__sro_n1316;
wire CLOCK_slo__sro_n1317;
wire CLOCK_slo__sro_n1318;
wire CLOCK_slo__sro_n1319;


INV_X1 i_36 (.ZN (n_34), .A (Multiplier[30]));
INV_X1 i_35 (.ZN (n_33), .A (p_0[30]));
INV_X1 i_34 (.ZN (n_32), .A (n_30));
OAI33_X1 i_33 (.ZN (n_31), .A1 (n_34), .A2 (p_0[30]), .A3 (n_32), .B1 (n_30), .B2 (n_33), .B3 (Multiplier[30]));
XOR2_X1 i_32 (.Z (p_1[31]), .A (Multiplier[31]), .B (n_31));
OAI22_X1 i_31 (.ZN (n_0), .A1 (n_34), .A2 (p_0[30]), .B1 (Multiplier[30]), .B2 (n_33));
XNOR2_X1 i_0 (.ZN (p_1[30]), .A (n_32), .B (n_0));
INV_X1 slo__sro_c21 (.ZN (slo__sro_n82), .A (slo__n168));
XNOR2_X1 CLOCK_slo__sro_c1044 (.ZN (p_1[15]), .A (n_15), .B (CLOCK_slo__sro_n1218));
INV_X1 slo__sro_c647 (.ZN (slo__sro_n763), .A (slo__sro_n778));
FA_X1 i_27 (.CO (n_27), .S (p_1[26]), .A (Multiplier[26]), .B (p_0[26]), .CI (n_26));
FA_X1 i_26 (.CO (n_26), .S (p_1[25]), .A (Multiplier[25]), .B (p_0[25]), .CI (n_25));
FA_X1 i_25 (.CO (n_25), .S (p_1[24]), .A (Multiplier[24]), .B (p_0[24]), .CI (n_24));
FA_X1 i_24 (.CO (n_24), .S (p_1[23]), .A (Multiplier[23]), .B (p_0[23]), .CI (n_23));
FA_X1 i_23 (.CO (n_23), .S (p_1[22]), .A (Multiplier[22]), .B (p_0[22]), .CI (n_22));
FA_X1 i_22 (.CO (n_22), .S (p_1[21]), .A (Multiplier[21]), .B (p_0[21]), .CI (n_21));
INV_X1 slo__sro_c663 (.ZN (slo__sro_n781), .A (n_19));
INV_X1 slo__sro_c698 (.ZN (slo__sro_n831), .A (n_4));
FA_X1 i_19 (.CO (n_19), .S (p_1[18]), .A (Multiplier[18]), .B (p_0[18]), .CI (n_18));
FA_X1 i_18 (.CO (n_18), .S (p_1[17]), .A (Multiplier[17]), .B (p_0[17]), .CI (slo__sro_n919));
NAND2_X2 CLOCK_slo__sro_c1030 (.ZN (slo__sro_n856), .A1 (n_8), .A2 (CLOCK_slo__sro_n1208));
INV_X1 CLOCK_slo__sro_c1212 (.ZN (CLOCK_slo__sro_n1405), .A (n_13));
NOR2_X1 CLOCK_slo__sro_c1214 (.ZN (CLOCK_slo__sro_n1403), .A1 (p_0[13]), .A2 (Multiplier[13]));
FA_X1 i_13 (.CO (n_13), .S (p_1[12]), .A (Multiplier[12]), .B (p_0[12]), .CI (n_12));
FA_X1 i_12 (.CO (n_12), .S (p_1[11]), .A (Multiplier[11]), .B (p_0[11]), .CI (CLOCK_slo__sro_n1316));
FA_X1 i_10 (.CO (n_10), .S (p_1[9]), .A (Multiplier[9]), .B (p_0[9]), .CI (n_9));
NAND2_X1 CLOCK_slo__sro_c1002 (.ZN (CLOCK_slo__sro_n1187), .A1 (p_0[3]), .A2 (Multiplier[3]));
FA_X1 i_8 (.CO (n_8), .S (p_1[7]), .A (Multiplier[7]), .B (p_0[7]), .CI (slo__sro_n79));
NAND2_X1 slo__sro_c35 (.ZN (slo__sro_n99), .A1 (p_0[1]), .A2 (Multiplier[1]));
NAND2_X1 slo__sro_c65 (.ZN (slo__sro_n129), .A1 (slo__sro_n96), .A2 (Multiplier[2]));
XNOR2_X2 slo__mro_c712 (.ZN (slo__mro_n844), .A (n_1), .B (Multiplier[1]));
INV_X1 CLOCK_slo__sro_c1039 (.ZN (CLOCK_slo__sro_n1222), .A (n_15));
INV_X1 slo__sro_c633 (.ZN (slo__sro_n748), .A (n_27));
INV_X1 slo__sro_c51 (.ZN (slo__sro_n117), .A (slo__sro_n828));
NAND2_X1 slo__sro_c150 (.ZN (slo__sro_n216), .A1 (p_0[28]), .A2 (Multiplier[28]));
INV_X1 slo__sro_c7 (.ZN (slo__sro_n66), .A (n_29));
NAND2_X1 slo__sro_c8 (.ZN (slo__sro_n65), .A1 (p_0[29]), .A2 (Multiplier[29]));
NOR2_X1 slo__sro_c9 (.ZN (slo__sro_n64), .A1 (p_0[29]), .A2 (Multiplier[29]));
OAI21_X1 slo__sro_c10 (.ZN (n_30), .A (slo__sro_n65), .B1 (slo__sro_n66), .B2 (slo__sro_n64));
XNOR2_X1 slo__sro_c11 (.ZN (slo__sro_n63), .A (p_0[29]), .B (Multiplier[29]));
XNOR2_X1 slo__sro_c12 (.ZN (p_1[29]), .A (n_29), .B (slo__sro_n63));
NAND2_X1 slo__sro_c22 (.ZN (slo__sro_n81), .A1 (p_0[6]), .A2 (Multiplier[6]));
NOR2_X1 slo__sro_c23 (.ZN (slo__sro_n80), .A1 (p_0[6]), .A2 (Multiplier[6]));
OAI21_X1 slo__sro_c24 (.ZN (slo__sro_n79), .A (slo__sro_n81), .B1 (slo__sro_n82), .B2 (slo__sro_n80));
XNOR2_X2 slo__sro_c25 (.ZN (slo__sro_n78), .A (p_0[6]), .B (Multiplier[6]));
XNOR2_X2 slo__sro_c26 (.ZN (p_1[6]), .A (slo__sro_n78), .B (n_6));
NAND2_X2 slo__sro_c36 (.ZN (slo__sro_n98), .A1 (n_1), .A2 (Multiplier[1]));
NAND2_X4 slo__sro_c37 (.ZN (slo__sro_n97), .A1 (p_0[1]), .A2 (n_1));
NAND3_X2 slo__sro_c38 (.ZN (slo__sro_n96), .A1 (slo__sro_n99), .A2 (slo__sro_n97), .A3 (slo__sro_n98));
NAND2_X1 slo__sro_c720 (.ZN (slo__sro_n857), .A1 (p_0[8]), .A2 (Multiplier[8]));
NAND2_X1 slo__sro_c634 (.ZN (slo__sro_n747), .A1 (p_0[27]), .A2 (Multiplier[27]));
NAND2_X1 slo__sro_c52 (.ZN (slo__sro_n116), .A1 (p_0[5]), .A2 (Multiplier[5]));
NOR2_X1 slo__sro_c53 (.ZN (slo__sro_n115), .A1 (p_0[5]), .A2 (Multiplier[5]));
OAI21_X1 slo__sro_c54 (.ZN (n_6), .A (slo__sro_n116), .B1 (slo__sro_n117), .B2 (slo__sro_n115));
XNOR2_X1 slo__sro_c55 (.ZN (slo__sro_n114), .A (p_0[5]), .B (Multiplier[5]));
XNOR2_X1 slo__sro_c56 (.ZN (p_1[5]), .A (slo__sro_n828), .B (slo__sro_n114));
OAI21_X1 slo__sro_c66 (.ZN (slo__sro_n128), .A (p_0[2]), .B1 (slo__sro_n96), .B2 (Multiplier[2]));
NAND2_X1 slo__sro_c67 (.ZN (n_3), .A1 (slo__sro_n128), .A2 (slo__sro_n129));
XNOR2_X1 slo__sro_c68 (.ZN (slo__sro_n127), .A (p_0[2]), .B (Multiplier[2]));
XNOR2_X2 slo__sro_c69 (.ZN (p_1[2]), .A (slo__sro_n127), .B (slo__sro_n96));
INV_X1 slo__sro_c149 (.ZN (slo__sro_n217), .A (n_28));
OAI21_X1 slo__c106 (.ZN (slo__n168), .A (slo__sro_n116), .B1 (slo__sro_n117), .B2 (slo__sro_n115));
INV_X1 slo__sro_c86 (.ZN (slo__sro_n148), .A (Multiplier[0]));
NAND2_X4 slo__sro_c87 (.ZN (slo__sro_n147), .A1 (p_0[0]), .A2 (Multiplier[0]));
INV_X4 slo__sro_c88 (.ZN (n_1), .A (slo__sro_n147));
XNOR2_X1 slo__sro_c89 (.ZN (p_1[0]), .A (opt_ipoPP_3), .B (slo__sro_n148));
NOR2_X1 slo__sro_c151 (.ZN (slo__sro_n215), .A1 (p_0[28]), .A2 (Multiplier[28]));
OAI21_X1 slo__sro_c152 (.ZN (n_29), .A (slo__sro_n216), .B1 (slo__sro_n217), .B2 (slo__sro_n215));
XNOR2_X1 slo__sro_c153 (.ZN (slo__sro_n214), .A (p_0[28]), .B (Multiplier[28]));
XNOR2_X1 slo__sro_c154 (.ZN (p_1[28]), .A (n_28), .B (slo__sro_n214));
NOR2_X1 slo__sro_c635 (.ZN (slo__sro_n746), .A1 (p_0[27]), .A2 (Multiplier[27]));
OAI21_X1 slo__sro_c636 (.ZN (n_28), .A (slo__sro_n747), .B1 (slo__sro_n748), .B2 (slo__sro_n746));
XNOR2_X1 slo__sro_c637 (.ZN (slo__sro_n745), .A (p_0[27]), .B (Multiplier[27]));
XNOR2_X1 slo__sro_c638 (.ZN (p_1[27]), .A (n_27), .B (slo__sro_n745));
NAND2_X1 slo__sro_c648 (.ZN (slo__sro_n762), .A1 (p_0[20]), .A2 (Multiplier[20]));
NOR2_X1 slo__sro_c649 (.ZN (slo__sro_n761), .A1 (p_0[20]), .A2 (Multiplier[20]));
OAI21_X1 slo__sro_c650 (.ZN (n_21), .A (slo__sro_n762), .B1 (slo__sro_n763), .B2 (slo__sro_n761));
XNOR2_X1 slo__sro_c651 (.ZN (slo__sro_n760), .A (p_0[20]), .B (Multiplier[20]));
XNOR2_X1 slo__sro_c652 (.ZN (p_1[20]), .A (slo__sro_n778), .B (slo__sro_n760));
NAND2_X1 slo__sro_c664 (.ZN (slo__sro_n780), .A1 (p_0[19]), .A2 (Multiplier[19]));
NOR2_X1 slo__sro_c665 (.ZN (slo__sro_n779), .A1 (p_0[19]), .A2 (Multiplier[19]));
OAI21_X1 slo__sro_c666 (.ZN (slo__sro_n778), .A (slo__sro_n780), .B1 (slo__sro_n781), .B2 (slo__sro_n779));
XNOR2_X1 slo__sro_c667 (.ZN (slo__sro_n777), .A (p_0[19]), .B (Multiplier[19]));
XNOR2_X1 slo__sro_c668 (.ZN (p_1[19]), .A (n_19), .B (slo__sro_n777));
NAND2_X1 slo__sro_c699 (.ZN (slo__sro_n830), .A1 (p_0[4]), .A2 (Multiplier[4]));
NOR2_X1 slo__sro_c700 (.ZN (slo__sro_n829), .A1 (p_0[4]), .A2 (Multiplier[4]));
OAI21_X2 slo__sro_c701 (.ZN (slo__sro_n828), .A (slo__sro_n830), .B1 (slo__sro_n831), .B2 (slo__sro_n829));
XNOR2_X1 slo__sro_c702 (.ZN (slo__sro_n827), .A (p_0[4]), .B (Multiplier[4]));
XNOR2_X1 slo__sro_c703 (.ZN (p_1[4]), .A (slo__sro_n827), .B (n_4));
XNOR2_X2 slo__mro_c713 (.ZN (p_1[1]), .A (slo__mro_n844), .B (p_0[1]));
NAND2_X2 slo__sro_c722 (.ZN (n_9), .A1 (slo__sro_n856), .A2 (slo__sro_n857));
XNOR2_X1 slo__sro_c723 (.ZN (slo__sro_n855), .A (p_0[8]), .B (Multiplier[8]));
XNOR2_X1 slo__sro_c724 (.ZN (p_1[8]), .A (slo__sro_n855), .B (n_8));
OAI21_X1 CLOCK_slo__sro_c1003 (.ZN (CLOCK_slo__sro_n1186), .A (n_3), .B1 (p_0[3]), .B2 (Multiplier[3]));
NAND2_X2 CLOCK_slo__sro_c1004 (.ZN (n_4), .A1 (CLOCK_slo__sro_n1186), .A2 (CLOCK_slo__sro_n1187));
XNOR2_X1 CLOCK_slo__sro_c1005 (.ZN (CLOCK_slo__sro_n1185), .A (p_0[3]), .B (Multiplier[3]));
XNOR2_X1 CLOCK_slo__sro_c1006 (.ZN (p_1[3]), .A (CLOCK_slo__sro_n1185), .B (n_3));
NAND2_X1 CLOCK_slo__sro_c1040 (.ZN (CLOCK_slo__sro_n1221), .A1 (Multiplier[15]), .A2 (p_0[15]));
NOR2_X1 CLOCK_slo__sro_c1041 (.ZN (CLOCK_slo__sro_n1220), .A1 (p_0[15]), .A2 (Multiplier[15]));
OAI21_X1 CLOCK_slo__sro_c1042 (.ZN (CLOCK_slo__sro_n1219), .A (CLOCK_slo__sro_n1221)
    , .B1 (CLOCK_slo__sro_n1222), .B2 (CLOCK_slo__sro_n1220));
XNOR2_X1 CLOCK_slo__sro_c1043 (.ZN (CLOCK_slo__sro_n1218), .A (p_0[15]), .B (Multiplier[15]));
INV_X1 CLOCK_slo__sro_c1027 (.ZN (CLOCK_slo__sro_n1210), .A (p_0[8]));
INV_X1 CLOCK_slo__sro_c1028 (.ZN (CLOCK_slo__sro_n1209), .A (Multiplier[8]));
NAND2_X1 CLOCK_slo__sro_c1029 (.ZN (CLOCK_slo__sro_n1208), .A1 (CLOCK_slo__sro_n1210), .A2 (CLOCK_slo__sro_n1209));
INV_X1 slo__sro_c782 (.ZN (slo__sro_n922), .A (CLOCK_slo__sro_n1219));
NAND2_X1 slo__sro_c783 (.ZN (slo__sro_n921), .A1 (Multiplier[16]), .A2 (p_0[16]));
NOR2_X1 slo__sro_c784 (.ZN (slo__sro_n920), .A1 (p_0[16]), .A2 (Multiplier[16]));
OAI21_X1 slo__sro_c785 (.ZN (slo__sro_n919), .A (slo__sro_n921), .B1 (slo__sro_n922), .B2 (slo__sro_n920));
XNOR2_X1 slo__sro_c786 (.ZN (slo__sro_n918), .A (p_0[16]), .B (Multiplier[16]));
XNOR2_X1 slo__sro_c787 (.ZN (p_1[16]), .A (CLOCK_slo__sro_n1219), .B (slo__sro_n918));
NAND2_X1 CLOCK_slo__sro_c1213 (.ZN (CLOCK_slo__sro_n1404), .A1 (p_0[13]), .A2 (Multiplier[13]));
NAND2_X1 CLOCK_slo__sro_c1073 (.ZN (CLOCK_slo__sro_n1258), .A1 (Multiplier[14]), .A2 (p_0[14]));
OR2_X1 CLOCK_slo__sro_c1074 (.ZN (CLOCK_slo__sro_n1257), .A1 (p_0[14]), .A2 (Multiplier[14]));
NAND2_X1 CLOCK_slo__sro_c1075 (.ZN (CLOCK_slo__sro_n1256), .A1 (CLOCK_slo__sro_n1402), .A2 (CLOCK_slo__sro_n1257));
NAND2_X1 CLOCK_slo__sro_c1076 (.ZN (n_15), .A1 (CLOCK_slo__sro_n1256), .A2 (CLOCK_slo__sro_n1258));
XNOR2_X1 CLOCK_slo__sro_c1077 (.ZN (CLOCK_slo__sro_n1255), .A (p_0[14]), .B (Multiplier[14]));
XNOR2_X1 CLOCK_slo__sro_c1078 (.ZN (p_1[14]), .A (CLOCK_slo__sro_n1402), .B (CLOCK_slo__sro_n1255));
OAI21_X1 CLOCK_slo__sro_c1215 (.ZN (CLOCK_slo__sro_n1402), .A (CLOCK_slo__sro_n1404)
    , .B1 (CLOCK_slo__sro_n1405), .B2 (CLOCK_slo__sro_n1403));
XNOR2_X1 CLOCK_slo__sro_c1216 (.ZN (CLOCK_slo__sro_n1401), .A (p_0[13]), .B (Multiplier[13]));
XNOR2_X1 CLOCK_slo__sro_c1217 (.ZN (p_1[13]), .A (n_13), .B (CLOCK_slo__sro_n1401));
INV_X2 CLOCK_slo__sro_c1132 (.ZN (CLOCK_slo__sro_n1319), .A (n_10));
NAND2_X1 CLOCK_slo__sro_c1133 (.ZN (CLOCK_slo__sro_n1318), .A1 (p_0[10]), .A2 (Multiplier[10]));
NOR2_X1 CLOCK_slo__sro_c1134 (.ZN (CLOCK_slo__sro_n1317), .A1 (p_0[10]), .A2 (Multiplier[10]));
OAI21_X2 CLOCK_slo__sro_c1135 (.ZN (CLOCK_slo__sro_n1316), .A (CLOCK_slo__sro_n1318)
    , .B1 (CLOCK_slo__sro_n1319), .B2 (CLOCK_slo__sro_n1317));
XNOR2_X1 CLOCK_slo__sro_c1136 (.ZN (CLOCK_slo__sro_n1315), .A (p_0[10]), .B (Multiplier[10]));
XNOR2_X1 CLOCK_slo__sro_c1137 (.ZN (p_1[10]), .A (n_10), .B (CLOCK_slo__sro_n1315));

endmodule //datapath__0_101

module datapath__0_96 (Multiplier, p_0, p_1);

output [31:0] p_1;
input [31:0] Multiplier;
input [31:0] p_0;
wire CLOCK_slo__sro_n1095;
wire slo__sro_n564;
wire slo__sro_n229;
wire n_1;
wire n_2;
wire n_4;
wire n_7;
wire n_8;
wire n_9;
wire n_11;
wire n_12;
wire n_13;
wire n_14;
wire n_15;
wire n_16;
wire n_17;
wire n_19;
wire n_20;
wire n_21;
wire n_23;
wire n_24;
wire n_25;
wire n_26;
wire n_28;
wire n_29;
wire n_30;
wire n_31;
wire slo__sro_n119;
wire slo__sro_n120;
wire slo__sro_n121;
wire slo__sro_n122;
wire slo__sro_n136;
wire slo__sro_n137;
wire slo__sro_n138;
wire slo__sro_n139;
wire slo__sro_n149;
wire slo__sro_n150;
wire slo__sro_n151;
wire slo__sro_n152;
wire slo__sro_n162;
wire slo__sro_n163;
wire slo__sro_n165;
wire slo__sro_n166;
wire slo__sro_n181;
wire slo__sro_n183;
wire slo__sro_n197;
wire slo__sro_n198;
wire slo__sro_n199;
wire slo__sro_n228;
wire slo__sro_n216;
wire slo__sro_n217;
wire slo__sro_n230;
wire slo__sro_n231;
wire slo__sro_n232;
wire slo__sro_n247;
wire slo__sro_n248;
wire slo__sro_n249;
wire slo__sro_n250;
wire slo__sro_n251;
wire slo__sro_n252;
wire slo__sro_n266;
wire slo__sro_n267;
wire slo__sro_n268;
wire slo__sro_n565;
wire slo__sro_n566;
wire opt_ipo_n513;
wire slo__sro_n567;
wire opt_ipo_n523;
wire slo__sro_n568;
wire slo__sro_n598;
wire slo__sro_n599;
wire slo__sro_n600;
wire slo__sro_n601;
wire slo__sro_n602;
wire slo__mro_n674;
wire CLOCK_slo__sro_n1105;
wire CLOCK_slo__sro_n1092;
wire CLOCK_slo__sro_n1093;
wire slo__n794;
wire CLOCK_slo__sro_n1094;
wire CLOCK_slo__sro_n1106;
wire CLOCK_slo__sro_n1107;
wire CLOCK_slo__sro_n1347;
wire CLOCK_slo__sro_n1226;
wire CLOCK_slo__sro_n1227;
wire CLOCK_slo__sro_n1228;
wire CLOCK_slo__sro_n1229;
wire CLOCK_slo__sro_n1230;
wire CLOCK_slo__sro_n1254;
wire CLOCK_slo__sro_n1255;
wire CLOCK_slo__sro_n1256;
wire CLOCK_slo__sro_n1257;
wire CLOCK_slo__sro_n1258;
wire CLOCK_slo__sro_n1348;
wire CLOCK_slo__sro_n1349;
wire CLOCK_slo__sro_n1350;
wire CLOCK_slo__sro_n1351;
wire CLOCK_slo__sro_n1513;


XNOR2_X1 i_32 (.ZN (p_1[31]), .A (n_31), .B (n_30));
XNOR2_X1 i_31 (.ZN (n_31), .A (Multiplier[31]), .B (p_0[31]));
FA_X1 i_30 (.CO (n_30), .S (p_1[30]), .A (Multiplier[30]), .B (p_0[30]), .CI (n_29));
NAND2_X1 slo__sro_c19 (.ZN (slo__sro_n139), .A1 (Multiplier[28]), .A2 (p_0[28]));
INV_X2 slo__sro_c33 (.ZN (slo__sro_n152), .A (n_12));
INV_X1 CLOCK_slo__sro_c964 (.ZN (CLOCK_slo__sro_n1258), .A (n_21));
FA_X1 i_26 (.CO (n_26), .S (p_1[26]), .A (Multiplier[26]), .B (p_0[26]), .CI (n_25));
FA_X1 i_25 (.CO (n_25), .S (p_1[25]), .A (Multiplier[25]), .B (p_0[25]), .CI (n_24));
FA_X1 i_24 (.CO (n_24), .S (p_1[24]), .A (Multiplier[24]), .B (p_0[24]), .CI (n_23));
FA_X1 i_23 (.CO (n_23), .S (p_1[23]), .A (Multiplier[23]), .B (p_0[23]), .CI (CLOCK_slo__sro_n1255));
INV_X2 CLOCK_slo__sro_c1057 (.ZN (CLOCK_slo__sro_n1351), .A (n_17));
FA_X1 i_21 (.CO (n_21), .S (p_1[21]), .A (Multiplier[21]), .B (p_0[21]), .CI (n_20));
FA_X1 i_20 (.CO (n_20), .S (p_1[20]), .A (Multiplier[20]), .B (p_0[20]), .CI (n_19));
FA_X1 i_19 (.CO (n_19), .S (p_1[19]), .A (Multiplier[19]), .B (p_0[19]), .CI (CLOCK_slo__sro_n1348));
FA_X1 i_17 (.CO (n_17), .S (p_1[17]), .A (Multiplier[17]), .B (p_0[17]), .CI (n_16));
FA_X1 i_16 (.CO (n_16), .S (p_1[16]), .A (Multiplier[16]), .B (p_0[16]), .CI (n_15));
FA_X1 i_15 (.CO (n_15), .S (p_1[15]), .A (Multiplier[15]), .B (p_0[15]), .CI (n_14));
FA_X1 i_14 (.CO (n_14), .S (p_1[14]), .A (Multiplier[14]), .B (p_0[14]), .CI (n_13));
INV_X4 slo__sro_c47 (.ZN (slo__sro_n166), .A (n_2));
INV_X2 slo__sro_c434 (.ZN (slo__sro_n602), .A (n_9));
NOR2_X1 CLOCK_slo__sro_c1059 (.ZN (CLOCK_slo__sro_n1349), .A1 (p_0[18]), .A2 (Multiplier[18]));
XNOR2_X1 CLOCK_slo__sro_c811 (.ZN (p_1[9]), .A (n_8), .B (CLOCK_slo__sro_n1092));
NAND2_X1 CLOCK_slo__sro_c820 (.ZN (CLOCK_slo__sro_n1107), .A1 (Multiplier[11]), .A2 (p_0[11]));
FA_X1 i_8 (.CO (n_8), .S (p_1[8]), .A (Multiplier[8]), .B (p_0[8]), .CI (n_7));
FA_X1 i_7 (.CO (n_7), .S (p_1[7]), .A (Multiplier[7]), .B (p_0[7]), .CI (slo__sro_n229));
NAND2_X1 slo__sro_c127 (.ZN (slo__sro_n252), .A1 (p_0[5]), .A2 (Multiplier[5]));
NAND2_X2 slo__sro_c143 (.ZN (slo__sro_n268), .A1 (slo__sro_n163), .A2 (Multiplier[4]));
NOR2_X1 slo__sro_c411 (.ZN (slo__sro_n567), .A1 (p_0[12]), .A2 (Multiplier[12]));
NAND2_X2 slo__sro_c63 (.ZN (slo__sro_n183), .A1 (n_1), .A2 (Multiplier[2]));
NAND2_X4 slo__sro_c78 (.ZN (slo__sro_n199), .A1 (opt_ipo_n513), .A2 (Multiplier[1]));
INV_X2 slo__sro_c111 (.ZN (slo__sro_n232), .A (slo__sro_n248));
XNOR2_X2 slo__sro_c115 (.ZN (slo__sro_n228), .A (p_0[6]), .B (Multiplier[6]));
INV_X1 slo__sro_c3 (.ZN (slo__sro_n122), .A (n_28));
NAND2_X1 slo__sro_c4 (.ZN (slo__sro_n121), .A1 (Multiplier[29]), .A2 (p_0[29]));
NOR2_X1 slo__sro_c5 (.ZN (slo__sro_n120), .A1 (p_0[29]), .A2 (Multiplier[29]));
OAI21_X1 slo__sro_c6 (.ZN (n_29), .A (slo__sro_n121), .B1 (slo__sro_n122), .B2 (slo__sro_n120));
XNOR2_X1 slo__sro_c7 (.ZN (slo__sro_n119), .A (p_0[29]), .B (Multiplier[29]));
XNOR2_X1 slo__sro_c8 (.ZN (p_1[29]), .A (n_28), .B (slo__sro_n119));
OR2_X1 slo__sro_c20 (.ZN (slo__sro_n138), .A1 (p_0[28]), .A2 (Multiplier[28]));
NAND2_X4 slo__sro_c21 (.ZN (slo__sro_n137), .A1 (CLOCK_slo__sro_n1227), .A2 (slo__sro_n138));
NAND2_X2 slo__sro_c22 (.ZN (n_28), .A1 (slo__sro_n137), .A2 (slo__sro_n139));
XNOR2_X1 slo__sro_c23 (.ZN (slo__sro_n136), .A (Multiplier[28]), .B (p_0[28]));
XNOR2_X1 slo__sro_c24 (.ZN (p_1[28]), .A (CLOCK_slo__sro_n1227), .B (slo__sro_n136));
NAND2_X1 slo__sro_c34 (.ZN (slo__sro_n151), .A1 (Multiplier[13]), .A2 (p_0[13]));
NOR2_X1 slo__sro_c35 (.ZN (slo__sro_n150), .A1 (p_0[13]), .A2 (Multiplier[13]));
OAI21_X2 slo__sro_c36 (.ZN (n_13), .A (slo__sro_n151), .B1 (slo__sro_n152), .B2 (slo__sro_n150));
XNOR2_X1 slo__sro_c37 (.ZN (slo__sro_n149), .A (Multiplier[13]), .B (p_0[13]));
XNOR2_X1 slo__sro_c38 (.ZN (p_1[13]), .A (n_12), .B (slo__sro_n149));
NAND2_X2 slo__sro_c48 (.ZN (slo__sro_n165), .A1 (p_0[3]), .A2 (Multiplier[3]));
INV_X2 CLOCK_slo__sro_c806 (.ZN (CLOCK_slo__sro_n1095), .A (n_8));
OAI21_X4 slo__sro_c50 (.ZN (slo__sro_n163), .A (slo__sro_n165), .B1 (slo__sro_n166), .B2 (slo__mro_n674));
XNOR2_X2 slo__sro_c51 (.ZN (slo__sro_n162), .A (p_0[3]), .B (Multiplier[3]));
XNOR2_X2 slo__sro_c52 (.ZN (p_1[3]), .A (slo__sro_n162), .B (n_2));
XNOR2_X2 slo__sro_c66 (.ZN (slo__sro_n181), .A (p_0[2]), .B (Multiplier[2]));
XNOR2_X2 slo__sro_c67 (.ZN (p_1[2]), .A (slo__sro_n181), .B (n_1));
OAI21_X4 slo__sro_c79 (.ZN (slo__sro_n198), .A (p_0[1]), .B1 (opt_ipo_n513), .B2 (Multiplier[1]));
NAND2_X2 slo__sro_c80 (.ZN (n_1), .A1 (slo__sro_n198), .A2 (slo__sro_n199));
XNOR2_X2 slo__sro_c81 (.ZN (slo__sro_n197), .A (p_0[1]), .B (Multiplier[1]));
XNOR2_X2 slo__sro_c82 (.ZN (p_1[1]), .A (slo__sro_n197), .B (opt_ipo_n513));
NAND2_X1 slo__sro_c112 (.ZN (slo__sro_n231), .A1 (Multiplier[6]), .A2 (p_0[6]));
NOR2_X2 slo__sro_c113 (.ZN (slo__sro_n230), .A1 (p_0[6]), .A2 (Multiplier[6]));
OAI21_X2 slo__sro_c114 (.ZN (slo__sro_n229), .A (slo__sro_n231), .B1 (slo__sro_n232), .B2 (slo__sro_n230));
INV_X1 slo__sro_c101 (.ZN (slo__sro_n217), .A (Multiplier[0]));
NAND2_X4 slo__sro_c102 (.ZN (slo__sro_n216), .A1 (p_0[0]), .A2 (Multiplier[0]));
NAND2_X1 slo__sro_c410 (.ZN (slo__sro_n568), .A1 (Multiplier[12]), .A2 (p_0[12]));
XNOR2_X1 slo__sro_c104 (.ZN (p_1[0]), .A (opt_ipo_n523), .B (slo__sro_n217));
XNOR2_X1 slo__sro_c116 (.ZN (p_1[6]), .A (slo__sro_n228), .B (slo__sro_n248));
NOR2_X1 slo__sro_c128 (.ZN (slo__sro_n251), .A1 (p_0[5]), .A2 (Multiplier[5]));
INV_X1 slo__sro_c129 (.ZN (slo__sro_n250), .A (slo__sro_n251));
NAND2_X2 slo__sro_c130 (.ZN (slo__sro_n249), .A1 (n_4), .A2 (slo__sro_n250));
NAND2_X2 slo__sro_c131 (.ZN (slo__sro_n248), .A1 (slo__sro_n249), .A2 (slo__sro_n252));
XNOR2_X1 slo__sro_c132 (.ZN (slo__sro_n247), .A (p_0[5]), .B (Multiplier[5]));
XNOR2_X1 slo__sro_c133 (.ZN (p_1[5]), .A (n_4), .B (slo__sro_n247));
AOI22_X4 slo__sro_c144 (.ZN (slo__sro_n267), .A1 (slo__sro_n163), .A2 (p_0[4]), .B1 (p_0[4]), .B2 (Multiplier[4]));
NAND2_X2 slo__sro_c145 (.ZN (n_4), .A1 (slo__sro_n267), .A2 (slo__sro_n268));
XNOR2_X2 slo__sro_c146 (.ZN (slo__sro_n266), .A (p_0[4]), .B (Multiplier[4]));
XNOR2_X2 slo__sro_c147 (.ZN (p_1[4]), .A (slo__sro_n163), .B (slo__sro_n266));
INV_X1 slo__sro_c412 (.ZN (slo__sro_n566), .A (slo__sro_n567));
NAND2_X2 slo__sro_c413 (.ZN (slo__sro_n565), .A1 (n_11), .A2 (slo__sro_n566));
INV_X4 opt_ipo_c382 (.ZN (opt_ipo_n513), .A (slo__sro_n216));
XNOR2_X1 slo__sro_c415 (.ZN (slo__sro_n564), .A (p_0[12]), .B (Multiplier[12]));
NAND2_X2 slo__sro_c414 (.ZN (n_12), .A1 (slo__sro_n565), .A2 (slo__sro_n568));
BUF_X1 opt_ipo_c392 (.Z (opt_ipo_n523), .A (p_0[0]));
XNOR2_X1 slo__sro_c416 (.ZN (p_1[12]), .A (n_11), .B (slo__sro_n564));
NAND2_X1 slo__sro_c435 (.ZN (slo__sro_n601), .A1 (Multiplier[10]), .A2 (p_0[10]));
NOR2_X2 slo__sro_c436 (.ZN (slo__sro_n600), .A1 (p_0[10]), .A2 (Multiplier[10]));
OAI21_X2 slo__sro_c437 (.ZN (slo__sro_n599), .A (slo__sro_n601), .B1 (slo__sro_n602), .B2 (slo__sro_n600));
XNOR2_X1 slo__sro_c438 (.ZN (slo__sro_n598), .A (p_0[10]), .B (Multiplier[10]));
XNOR2_X1 slo__sro_c439 (.ZN (p_1[10]), .A (n_9), .B (slo__sro_n598));
OAI21_X2 CLOCK_slo__sro_c821 (.ZN (CLOCK_slo__sro_n1106), .A (slo__sro_n599), .B1 (p_0[11]), .B2 (Multiplier[11]));
NOR2_X4 slo__mro_c506 (.ZN (slo__mro_n674), .A1 (p_0[3]), .A2 (Multiplier[3]));
NAND2_X1 CLOCK_slo__sro_c807 (.ZN (CLOCK_slo__sro_n1094), .A1 (p_0[9]), .A2 (Multiplier[9]));
NOR2_X2 CLOCK_slo__sro_c808 (.ZN (CLOCK_slo__sro_n1093), .A1 (p_0[9]), .A2 (Multiplier[9]));
OAI21_X2 CLOCK_slo__sro_c809 (.ZN (n_9), .A (CLOCK_slo__sro_n1094), .B1 (CLOCK_slo__sro_n1095), .B2 (CLOCK_slo__sro_n1093));
XNOR2_X1 CLOCK_slo__sro_c810 (.ZN (CLOCK_slo__sro_n1092), .A (p_0[9]), .B (Multiplier[9]));
NAND2_X4 slo__c597 (.ZN (slo__n794), .A1 (slo__sro_n198), .A2 (slo__sro_n199));
NAND2_X4 CLOCK_slo__sro_c822 (.ZN (n_11), .A1 (CLOCK_slo__sro_n1106), .A2 (CLOCK_slo__sro_n1107));
XNOR2_X1 CLOCK_slo__sro_c823 (.ZN (CLOCK_slo__sro_n1105), .A (p_0[11]), .B (Multiplier[11]));
XNOR2_X1 CLOCK_slo__sro_c824 (.ZN (p_1[11]), .A (CLOCK_slo__sro_n1105), .B (slo__sro_n599));
INV_X1 CLOCK_slo__sro_c946 (.ZN (CLOCK_slo__sro_n1230), .A (n_26));
NAND2_X1 CLOCK_slo__sro_c947 (.ZN (CLOCK_slo__sro_n1229), .A1 (p_0[27]), .A2 (Multiplier[27]));
NOR2_X1 CLOCK_slo__sro_c948 (.ZN (CLOCK_slo__sro_n1228), .A1 (Multiplier[27]), .A2 (p_0[27]));
OAI21_X2 CLOCK_slo__sro_c949 (.ZN (CLOCK_slo__sro_n1227), .A (CLOCK_slo__sro_n1229)
    , .B1 (CLOCK_slo__sro_n1230), .B2 (CLOCK_slo__sro_n1228));
XNOR2_X1 CLOCK_slo__sro_c950 (.ZN (CLOCK_slo__sro_n1226), .A (p_0[27]), .B (Multiplier[27]));
XNOR2_X1 CLOCK_slo__sro_c951 (.ZN (p_1[27]), .A (n_26), .B (CLOCK_slo__sro_n1226));
NAND2_X1 CLOCK_slo__sro_c965 (.ZN (CLOCK_slo__sro_n1257), .A1 (Multiplier[22]), .A2 (p_0[22]));
NOR2_X1 CLOCK_slo__sro_c966 (.ZN (CLOCK_slo__sro_n1256), .A1 (p_0[22]), .A2 (Multiplier[22]));
OAI21_X1 CLOCK_slo__sro_c967 (.ZN (CLOCK_slo__sro_n1255), .A (CLOCK_slo__sro_n1257)
    , .B1 (CLOCK_slo__sro_n1258), .B2 (CLOCK_slo__sro_n1256));
XNOR2_X1 CLOCK_slo__sro_c968 (.ZN (CLOCK_slo__sro_n1254), .A (p_0[22]), .B (Multiplier[22]));
XNOR2_X1 CLOCK_slo__sro_c969 (.ZN (p_1[22]), .A (n_21), .B (CLOCK_slo__sro_n1254));
NAND2_X1 CLOCK_slo__sro_c1058 (.ZN (CLOCK_slo__sro_n1350), .A1 (Multiplier[18]), .A2 (p_0[18]));
OAI21_X1 CLOCK_slo__sro_c1060 (.ZN (CLOCK_slo__sro_n1348), .A (CLOCK_slo__sro_n1350)
    , .B1 (CLOCK_slo__sro_n1351), .B2 (CLOCK_slo__sro_n1349));
XNOR2_X1 CLOCK_slo__sro_c1061 (.ZN (CLOCK_slo__sro_n1347), .A (p_0[18]), .B (Multiplier[18]));
XNOR2_X1 CLOCK_slo__sro_c1062 (.ZN (p_1[18]), .A (n_17), .B (CLOCK_slo__sro_n1347));
OAI21_X4 CLOCK_slo__sro_c1224 (.ZN (CLOCK_slo__sro_n1513), .A (p_0[2]), .B1 (slo__n794), .B2 (Multiplier[2]));
NAND2_X4 CLOCK_slo__mro_c1215 (.ZN (n_2), .A1 (slo__sro_n183), .A2 (CLOCK_slo__sro_n1513));

endmodule //datapath__0_96

module datapath (p_0_18_PP_1, p_0_18_PP_2, p_0_19_PP_1, p_0_24_PP_2, drc_ipoPP_0, 
    Multiplier, p_0);

output [31:0] p_0;
output p_0_18_PP_1;
output p_0_18_PP_2;
output p_0_19_PP_1;
output p_0_24_PP_2;
input [31:0] Multiplier;
input drc_ipoPP_0;
wire drc_ipo_n106;
wire drc_ipo_n108;
wire drc_ipo_n110;
wire drc_ipo_n112;
wire drc_ipo_n114;
wire drc_ipo_n116;
wire drc_ipo_n118;
wire drc_ipo_n120;
wire drc_ipo_n122;
wire drc_ipo_n124;
wire drc_ipo_n126;
wire drc_ipo_n128;
wire drc_ipo_n130;
wire drc_ipo_n132;
wire drc_ipo_n134;
wire drc_ipo_n136;
wire drc_ipo_n138;
wire drc_ipo_n140;
wire drc_ipo_n142;
wire drc_ipo_n144;
wire drc_ipo_n146;
wire drc_ipo_n148;
wire drc_ipo_n150;
wire slo__n469;
wire drc_ipo_n154;
wire slo__n408;
wire CLOCK_spc__n1636;
wire n_0;
wire CLOCK_opt_ipo_n1207;
wire n_28;
wire n_27;
wire n_26;
wire n_25;
wire n_24;
wire n_1;
wire n_23;
wire n_22;
wire n_21;
wire n_20;
wire n_19;
wire n_18;
wire n_2;
wire n_17;
wire n_16;
wire n_15;
wire n_14;
wire n_13;
wire n_12;
wire n_11;
wire n_9;
wire n_3;
wire n_10;
wire n_8;
wire n_7;
wire n_6;
wire n_5;
wire n_4;
wire n_34;
wire n_33;
wire n_32;
wire n_31;
wire sgo__n215;
wire sgo__n307;
wire sgo__n227;
wire sgo__n228;
wire sgo__n243;
wire sgo__n244;
wire sgo__n265;
wire sgo__n266;
wire slo__mro_n340;
wire slo__sro_n437;
wire slo__sro_n438;
wire slo__sro_n492;
wire slo__sro_n577;
wire slo__sro_n578;
wire CLOCK_spc__n1635;
wire slo__sro_n579;
wire slo__sro_n580;
wire opt_ipo_n743;
wire CLOCK_spc__n1634;

// WARNING . Detected multiport output net(s). Introducing ASSIGN statements.
// This may cause simulation/synthesis mismatches . 
assign p_0[24] = p_0_24_PP_2;
assign p_0[19] = p_0_19_PP_1;
assign p_0[18] = p_0_18_PP_2;
assign p_0_18_PP_1 = p_0_18_PP_2;

INV_X1 i_65 (.ZN (n_34), .A (Multiplier[27]));
INV_X1 i_64 (.ZN (n_33), .A (Multiplier[21]));
INV_X1 i_63 (.ZN (n_32), .A (Multiplier[14]));
INV_X1 i_62 (.ZN (n_31), .A (Multiplier[6]));
XNOR2_X2 slo__mro_c126 (.ZN (p_0[1]), .A (slo__mro_n340), .B (Multiplier[0]));
INV_X1 slo__sro_c225 (.ZN (slo__sro_n438), .A (Multiplier[4]));
NOR2_X2 i_59 (.ZN (n_28), .A1 (CLOCK_opt_ipo_n1207), .A2 (Multiplier[4]));
NOR3_X2 i_58 (.ZN (n_27), .A1 (CLOCK_opt_ipo_n1207), .A2 (Multiplier[4]), .A3 (Multiplier[5]));
NAND2_X1 i_57 (.ZN (n_26), .A1 (slo__sro_n577), .A2 (n_31));
OR2_X2 i_56 (.ZN (n_25), .A1 (n_26), .A2 (Multiplier[7]));
INV_X1 slo__sro_c262 (.ZN (slo__sro_n492), .A (Multiplier[3]));
OR2_X1 i_54 (.ZN (n_23), .A1 (n_24), .A2 (Multiplier[10]));
OR2_X1 i_53 (.ZN (n_22), .A1 (n_23), .A2 (drc_ipoPP_0));
NOR2_X1 i_52 (.ZN (n_21), .A1 (n_22), .A2 (Multiplier[12]));
NOR3_X2 i_51 (.ZN (n_20), .A1 (n_22), .A2 (Multiplier[12]), .A3 (Multiplier[13]));
NAND2_X1 i_50 (.ZN (n_19), .A1 (n_20), .A2 (n_32));
OR3_X1 i_49 (.ZN (n_18), .A1 (n_19), .A2 (Multiplier[15]), .A3 (Multiplier[16]));
OR2_X1 i_48 (.ZN (n_17), .A1 (n_18), .A2 (Multiplier[17]));
NOR2_X1 i_47 (.ZN (n_16), .A1 (n_17), .A2 (Multiplier[18]));
NOR3_X1 i_46 (.ZN (n_15), .A1 (n_17), .A2 (Multiplier[18]), .A3 (Multiplier[19]));
NOR4_X1 i_45 (.ZN (n_14), .A1 (n_17), .A2 (Multiplier[18]), .A3 (Multiplier[19]), .A4 (Multiplier[20]));
NAND2_X1 i_44 (.ZN (n_13), .A1 (CLOCK_spc__n1636), .A2 (n_33));
OR2_X1 i_43 (.ZN (n_12), .A1 (n_13), .A2 (Multiplier[22]));
NOR2_X1 i_42 (.ZN (n_11), .A1 (n_12), .A2 (Multiplier[23]));
INV_X1 i_41 (.ZN (n_10), .A (n_11));
OR3_X1 i_40 (.ZN (n_9), .A1 (n_10), .A2 (Multiplier[24]), .A3 (Multiplier[25]));
NOR2_X1 i_39 (.ZN (n_8), .A1 (n_9), .A2 (Multiplier[26]));
NAND2_X1 i_38 (.ZN (n_7), .A1 (n_8), .A2 (n_34));
NOR2_X1 i_37 (.ZN (n_6), .A1 (n_7), .A2 (Multiplier[28]));
NOR3_X1 i_36 (.ZN (n_5), .A1 (n_7), .A2 (Multiplier[28]), .A3 (Multiplier[29]));
NOR4_X1 i_35 (.ZN (n_4), .A1 (n_7), .A2 (Multiplier[28]), .A3 (Multiplier[29]), .A4 (Multiplier[30]));
XNOR2_X1 i_34 (.ZN (drc_ipo_n106), .A (Multiplier[31]), .B (n_4));
XNOR2_X2 i_33 (.ZN (p_0[30]), .A (Multiplier[30]), .B (n_5));
XNOR2_X1 i_32 (.ZN (drc_ipo_n108), .A (Multiplier[29]), .B (n_6));
XOR2_X2 i_31 (.Z (drc_ipo_n110), .A (Multiplier[28]), .B (n_7));
XNOR2_X2 i_30 (.ZN (drc_ipo_n112), .A (Multiplier[27]), .B (n_8));
XOR2_X2 i_29 (.Z (drc_ipo_n114), .A (Multiplier[26]), .B (n_9));
OAI21_X1 i_28 (.ZN (n_3), .A (Multiplier[25]), .B1 (n_10), .B2 (Multiplier[24]));
AND2_X1 i_27 (.ZN (sgo__n265), .A1 (n_9), .A2 (n_3));
XNOR2_X1 i_26 (.ZN (drc_ipo_n116), .A (Multiplier[24]), .B (n_11));
XOR2_X2 i_25 (.Z (drc_ipo_n118), .A (Multiplier[23]), .B (n_12));
XOR2_X1 i_24 (.Z (drc_ipo_n120), .A (Multiplier[22]), .B (n_13));
XNOR2_X2 i_23 (.ZN (drc_ipo_n122), .A (Multiplier[21]), .B (CLOCK_spc__n1635));
XNOR2_X1 i_22 (.ZN (drc_ipo_n124), .A (Multiplier[20]), .B (n_15));
XNOR2_X1 i_21 (.ZN (drc_ipo_n126), .A (Multiplier[19]), .B (n_16));
XOR2_X1 i_20 (.Z (drc_ipo_n128), .A (Multiplier[18]), .B (n_17));
XOR2_X1 i_19 (.Z (drc_ipo_n130), .A (Multiplier[17]), .B (n_18));
OAI21_X1 i_18 (.ZN (n_2), .A (Multiplier[16]), .B1 (n_19), .B2 (Multiplier[15]));
AND2_X1 i_17 (.ZN (sgo__n243), .A1 (n_18), .A2 (n_2));
XOR2_X1 i_16 (.Z (drc_ipo_n132), .A (Multiplier[15]), .B (n_19));
XNOR2_X2 i_15 (.ZN (drc_ipo_n134), .A (Multiplier[14]), .B (n_20));
XNOR2_X2 i_14 (.ZN (drc_ipo_n136), .A (Multiplier[13]), .B (n_21));
XOR2_X2 i_13 (.Z (drc_ipo_n138), .A (Multiplier[12]), .B (n_22));
XOR2_X2 i_12 (.Z (drc_ipo_n140), .A (Multiplier[11]), .B (n_23));
XOR2_X1 i_11 (.Z (drc_ipo_n142), .A (Multiplier[10]), .B (n_24));
OAI21_X1 i_10 (.ZN (n_1), .A (Multiplier[9]), .B1 (n_25), .B2 (Multiplier[8]));
AND2_X1 i_9 (.ZN (sgo__n227), .A1 (n_24), .A2 (n_1));
XOR2_X1 i_8 (.Z (drc_ipo_n144), .A (Multiplier[8]), .B (n_25));
XOR2_X1 i_7 (.Z (drc_ipo_n146), .A (Multiplier[7]), .B (n_26));
XNOR2_X1 i_6 (.ZN (drc_ipo_n148), .A (n_27), .B (Multiplier[6]));
XNOR2_X1 i_5 (.ZN (drc_ipo_n150), .A (n_28), .B (Multiplier[5]));
NOR3_X1 slo__c245 (.ZN (slo__n469), .A1 (n_25), .A2 (Multiplier[8]), .A3 (Multiplier[9]));
INV_X4 CLOCK_opt_ipo_c674 (.ZN (CLOCK_opt_ipo_n1207), .A (slo__n408));
OAI21_X1 i_2 (.ZN (n_0), .A (Multiplier[2]), .B1 (Multiplier[0]), .B2 (Multiplier[1]));
NOR3_X4 sgo__c109 (.ZN (sgo__n307), .A1 (Multiplier[0]), .A2 (Multiplier[1]), .A3 (Multiplier[2]));
NOR2_X4 slo__c188 (.ZN (slo__n408), .A1 (opt_ipo_n743), .A2 (Multiplier[3]));
BUF_X8 drc_ipo_c53 (.Z (p_0[31]), .A (drc_ipo_n106));
BUF_X2 drc_ipo_c54 (.Z (p_0[29]), .A (drc_ipo_n108));
BUF_X32 drc_ipo_c55 (.Z (p_0[28]), .A (drc_ipo_n110));
BUF_X32 drc_ipo_c56 (.Z (p_0[27]), .A (drc_ipo_n112));
BUF_X32 drc_ipo_c57 (.Z (p_0[26]), .A (drc_ipo_n114));
BUF_X4 drc_ipo_c58 (.Z (p_0_24_PP_2), .A (drc_ipo_n116));
BUF_X32 drc_ipo_c59 (.Z (p_0[23]), .A (drc_ipo_n118));
BUF_X8 drc_ipo_c60 (.Z (p_0[22]), .A (drc_ipo_n120));
BUF_X32 drc_ipo_c61 (.Z (p_0[21]), .A (drc_ipo_n122));
BUF_X8 drc_ipo_c62 (.Z (p_0[20]), .A (drc_ipo_n124));
BUF_X8 drc_ipo_c63 (.Z (p_0_19_PP_1), .A (drc_ipo_n126));
BUF_X4 drc_ipo_c64 (.Z (p_0_18_PP_2), .A (drc_ipo_n128));
BUF_X8 drc_ipo_c65 (.Z (p_0[17]), .A (drc_ipo_n130));
BUF_X8 drc_ipo_c66 (.Z (p_0[15]), .A (drc_ipo_n132));
BUF_X32 drc_ipo_c67 (.Z (p_0[14]), .A (drc_ipo_n134));
BUF_X32 drc_ipo_c68 (.Z (p_0[13]), .A (drc_ipo_n136));
BUF_X32 drc_ipo_c69 (.Z (p_0[12]), .A (drc_ipo_n138));
BUF_X32 drc_ipo_c70 (.Z (p_0[11]), .A (drc_ipo_n140));
BUF_X8 drc_ipo_c71 (.Z (p_0[10]), .A (drc_ipo_n142));
BUF_X8 drc_ipo_c72 (.Z (p_0[8]), .A (drc_ipo_n144));
BUF_X4 drc_ipo_c73 (.Z (p_0[7]), .A (drc_ipo_n146));
BUF_X4 drc_ipo_c74 (.Z (p_0[6]), .A (drc_ipo_n148));
BUF_X4 drc_ipo_c75 (.Z (p_0[5]), .A (drc_ipo_n150));
BUF_X4 drc_ipo_c76 (.Z (p_0[4]), .A (slo__sro_n437));
BUF_X4 drc_ipo_c77 (.Z (p_0[3]), .A (drc_ipo_n154));
INV_X2 opt_ipo_c447 (.ZN (opt_ipo_n743), .A (sgo__n307));
INV_X4 sgo__c80 (.ZN (p_0[2]), .A (sgo__n215));
INV_X1 sgo__c81 (.ZN (sgo__n228), .A (sgo__n227));
INV_X4 sgo__c82 (.ZN (p_0[9]), .A (sgo__n228));
INV_X2 sgo__c83 (.ZN (sgo__n244), .A (sgo__n243));
INV_X32 sgo__c84 (.ZN (p_0[16]), .A (sgo__n244));
INV_X1 sgo__c85 (.ZN (sgo__n266), .A (sgo__n265));
INV_X2 sgo__c86 (.ZN (p_0[25]), .A (sgo__n266));
INV_X2 slo__mro_c125 (.ZN (slo__mro_n340), .A (Multiplier[1]));
NAND2_X2 sgo__c100 (.ZN (sgo__n215), .A1 (opt_ipo_n743), .A2 (n_0));
INV_X1 CLOCK_spc__L1_c930 (.ZN (CLOCK_spc__n1634), .A (n_14));
XNOR2_X2 slo__sro_c226 (.ZN (slo__sro_n437), .A (CLOCK_opt_ipo_n1207), .B (slo__sro_n438));
INV_X1 slo__c247 (.ZN (n_24), .A (slo__n469));
XNOR2_X2 slo__sro_c263 (.ZN (drc_ipo_n154), .A (opt_ipo_n743), .B (slo__sro_n492));
INV_X1 slo__sro_c344 (.ZN (slo__sro_n580), .A (Multiplier[4]));
INV_X1 slo__sro_c345 (.ZN (slo__sro_n579), .A (Multiplier[5]));
NAND2_X1 slo__sro_c346 (.ZN (slo__sro_n578), .A1 (slo__sro_n579), .A2 (slo__sro_n580));
NOR2_X1 slo__sro_c347 (.ZN (slo__sro_n577), .A1 (CLOCK_opt_ipo_n1207), .A2 (slo__sro_n578));
INV_X1 CLOCK_spc__L2_c931 (.ZN (CLOCK_spc__n1635), .A (CLOCK_spc__n1634));
INV_X1 CLOCK_spc__L2_c932 (.ZN (CLOCK_spc__n1636), .A (CLOCK_spc__n1634));

endmodule //datapath

module BoothAlgorithmMultiplier (Multiplier_0_PP_0, drc_ipoPP_0, drc_ipoPP_1, drc_ipoPP_2, 
    drc_ipoPP_3, drc_ipoPP_4, drc_ipoPP_5, drc_ipoPP_6, drc_ipoPP_7, Multiplier_19_PP_2, 
    drc_ipoPP_3PP_0, drc_ipoPP_2PP_0, Multiplicand, Multiplier, Product);

output [63:0] Product;
input [31:0] Multiplicand;
input [31:0] Multiplier;
input Multiplier_0_PP_0;
input drc_ipoPP_0;
input drc_ipoPP_1;
input drc_ipoPP_2;
input drc_ipoPP_3;
input drc_ipoPP_4;
input drc_ipoPP_5;
input drc_ipoPP_6;
input drc_ipoPP_7;
input Multiplier_19_PP_2;
input drc_ipoPP_3PP_0;
input drc_ipoPP_2PP_0;
wire CLOCK_sgo__n46725;
wire opt_ipo_n43864;
wire slo__sro_n39796;
wire n_6_0;
wire n_6_1;
wire n_6_2;
wire n_6_3;
wire n_6_4;
wire n_6_5;
wire n_6_6;
wire n_6_7;
wire n_6_8;
wire n_6_9;
wire n_6_10;
wire n_6_11;
wire n_6_12;
wire n_6_13;
wire n_6_14;
wire n_6_15;
wire n_6_16;
wire n_6_17;
wire CLOCK_slo__mro_n62209;
wire n_6_19;
wire n_6_20;
wire n_6_21;
wire n_6_22;
wire n_6_23;
wire n_6_24;
wire n_6_25;
wire n_6_26;
wire n_6_27;
wire n_6_28;
wire n_6_29;
wire n_6_30;
wire n_6_31;
wire n_6_32;
wire n_6_33;
wire n_6_34;
wire n_6_35;
wire n_6_36;
wire n_6_37;
wire n_6_38;
wire n_6_39;
wire n_6_40;
wire n_6_41;
wire n_6_42;
wire n_6_43;
wire n_6_44;
wire n_6_45;
wire n_6_46;
wire n_6_47;
wire n_6_48;
wire n_6_49;
wire n_6_50;
wire n_6_51;
wire n_6_52;
wire n_6_53;
wire n_6_54;
wire n_6_55;
wire n_6_56;
wire n_6_57;
wire n_6_58;
wire n_6_59;
wire n_6_60;
wire n_6_61;
wire n_6_62;
wire n_6_63;
wire n_6_64;
wire n_6_65;
wire n_6_66;
wire n_6_67;
wire n_6_68;
wire n_6_69;
wire n_6_70;
wire n_6_71;
wire n_6_72;
wire n_6_73;
wire n_6_74;
wire n_6_75;
wire n_6_76;
wire n_6_77;
wire n_6_78;
wire n_6_79;
wire n_6_80;
wire n_6_81;
wire n_6_82;
wire n_6_83;
wire n_6_84;
wire n_6_85;
wire n_6_86;
wire n_6_87;
wire n_6_88;
wire n_6_89;
wire n_6_90;
wire n_6_91;
wire n_6_92;
wire n_6_93;
wire n_6_94;
wire n_6_95;
wire n_6_96;
wire n_6_97;
wire n_6_98;
wire n_6_99;
wire n_6_100;
wire n_6_101;
wire n_6_102;
wire n_6_103;
wire n_6_104;
wire n_6_105;
wire n_6_106;
wire n_6_107;
wire n_6_108;
wire n_6_109;
wire n_6_110;
wire n_6_111;
wire n_6_112;
wire n_6_113;
wire n_6_114;
wire n_6_115;
wire n_6_116;
wire n_6_117;
wire n_6_118;
wire n_6_119;
wire n_6_120;
wire n_6_121;
wire n_6_122;
wire n_6_123;
wire n_6_124;
wire n_6_125;
wire n_6_126;
wire n_6_127;
wire n_6_128;
wire n_6_129;
wire n_6_130;
wire n_6_131;
wire n_6_132;
wire n_6_133;
wire n_6_134;
wire n_6_135;
wire n_6_136;
wire n_6_137;
wire n_6_138;
wire n_6_139;
wire n_6_140;
wire n_6_141;
wire n_6_142;
wire n_6_143;
wire n_6_144;
wire n_6_145;
wire n_6_146;
wire n_6_147;
wire n_6_148;
wire n_6_149;
wire n_6_150;
wire n_6_151;
wire n_6_152;
wire n_6_153;
wire n_6_154;
wire n_6_155;
wire n_6_156;
wire n_6_157;
wire n_6_158;
wire n_6_159;
wire n_6_160;
wire n_6_161;
wire n_6_162;
wire n_6_163;
wire n_6_164;
wire n_6_165;
wire n_6_166;
wire n_6_167;
wire n_6_168;
wire n_6_169;
wire n_6_170;
wire n_6_171;
wire n_6_172;
wire n_6_173;
wire n_6_174;
wire n_6_175;
wire n_6_176;
wire n_6_177;
wire n_6_178;
wire n_6_179;
wire n_6_180;
wire n_6_181;
wire n_6_182;
wire n_6_183;
wire n_6_184;
wire n_6_185;
wire n_6_186;
wire n_6_187;
wire n_6_188;
wire n_6_189;
wire n_6_190;
wire n_6_191;
wire n_6_192;
wire n_6_193;
wire n_6_194;
wire n_6_195;
wire n_6_196;
wire n_6_197;
wire n_6_198;
wire n_6_199;
wire n_6_200;
wire n_6_201;
wire n_6_202;
wire n_6_203;
wire n_6_204;
wire n_6_205;
wire n_6_206;
wire n_6_207;
wire n_6_208;
wire n_6_209;
wire n_6_210;
wire n_6_211;
wire n_6_212;
wire n_6_213;
wire n_6_214;
wire n_6_215;
wire n_6_216;
wire n_6_217;
wire n_6_218;
wire n_6_219;
wire n_6_220;
wire n_6_221;
wire n_6_222;
wire n_6_223;
wire n_6_224;
wire n_6_225;
wire n_6_226;
wire n_6_227;
wire n_6_228;
wire n_6_229;
wire n_6_230;
wire n_6_231;
wire n_6_232;
wire n_6_233;
wire n_6_234;
wire n_6_235;
wire n_6_236;
wire n_6_237;
wire n_6_238;
wire n_6_239;
wire n_6_240;
wire n_6_241;
wire n_6_242;
wire n_6_243;
wire n_6_244;
wire n_6_245;
wire n_6_246;
wire n_6_247;
wire n_6_248;
wire n_6_249;
wire n_6_250;
wire n_6_251;
wire n_6_252;
wire n_6_253;
wire n_6_254;
wire n_6_255;
wire n_6_256;
wire n_6_257;
wire n_6_258;
wire n_6_259;
wire n_6_260;
wire n_6_261;
wire n_6_262;
wire n_6_263;
wire n_6_264;
wire n_6_265;
wire n_6_266;
wire n_6_267;
wire n_6_268;
wire n_6_269;
wire n_6_270;
wire n_6_271;
wire n_6_272;
wire n_6_273;
wire n_6_274;
wire n_6_275;
wire n_6_276;
wire n_6_277;
wire n_6_278;
wire n_6_279;
wire n_6_280;
wire n_6_281;
wire n_6_282;
wire n_6_283;
wire n_6_284;
wire n_6_285;
wire n_6_286;
wire n_6_287;
wire n_6_288;
wire n_6_289;
wire n_6_290;
wire n_6_291;
wire n_6_292;
wire n_6_293;
wire n_6_294;
wire n_6_295;
wire n_6_296;
wire n_6_297;
wire n_6_298;
wire n_6_299;
wire n_6_300;
wire n_6_301;
wire n_6_302;
wire n_6_303;
wire n_6_304;
wire n_6_305;
wire n_6_306;
wire n_6_307;
wire n_6_308;
wire n_6_309;
wire n_6_310;
wire n_6_311;
wire n_6_312;
wire n_6_313;
wire n_6_314;
wire n_6_315;
wire n_6_316;
wire n_6_317;
wire n_6_318;
wire n_6_319;
wire n_6_320;
wire n_6_321;
wire n_6_322;
wire n_6_323;
wire n_6_324;
wire n_6_325;
wire n_6_326;
wire n_6_327;
wire n_6_328;
wire n_6_329;
wire n_6_330;
wire n_6_331;
wire n_6_332;
wire n_6_333;
wire n_6_334;
wire n_6_335;
wire n_6_336;
wire n_6_337;
wire n_6_338;
wire n_6_339;
wire n_6_340;
wire n_6_341;
wire n_6_342;
wire n_6_343;
wire n_6_344;
wire n_6_345;
wire n_6_346;
wire n_6_347;
wire n_6_348;
wire n_6_349;
wire n_6_350;
wire n_6_351;
wire n_6_352;
wire n_6_353;
wire n_6_354;
wire n_6_355;
wire n_6_356;
wire n_6_357;
wire n_6_358;
wire n_6_359;
wire n_6_360;
wire n_6_361;
wire n_6_362;
wire n_6_363;
wire n_6_364;
wire n_6_365;
wire n_6_366;
wire n_6_367;
wire n_6_368;
wire n_6_369;
wire n_6_370;
wire n_6_371;
wire n_6_372;
wire n_6_373;
wire n_6_374;
wire n_6_375;
wire n_6_376;
wire n_6_377;
wire n_6_378;
wire n_6_379;
wire n_6_380;
wire n_6_381;
wire n_6_382;
wire n_6_383;
wire n_6_384;
wire n_6_385;
wire n_6_386;
wire n_6_387;
wire n_6_388;
wire n_6_389;
wire n_6_390;
wire n_6_391;
wire n_6_392;
wire n_6_393;
wire n_6_394;
wire n_6_395;
wire n_6_396;
wire n_6_397;
wire n_6_398;
wire n_6_399;
wire n_6_400;
wire n_6_401;
wire n_6_402;
wire n_6_403;
wire n_6_404;
wire n_6_405;
wire n_6_406;
wire n_6_407;
wire n_6_408;
wire n_6_409;
wire n_6_410;
wire n_6_411;
wire n_6_412;
wire n_6_413;
wire n_6_414;
wire n_6_415;
wire n_6_416;
wire n_6_417;
wire n_6_418;
wire n_6_419;
wire n_6_420;
wire n_6_421;
wire n_6_422;
wire n_6_423;
wire n_6_424;
wire n_6_425;
wire n_6_426;
wire n_6_427;
wire n_6_428;
wire n_6_429;
wire n_6_430;
wire n_6_431;
wire n_6_432;
wire n_6_433;
wire n_6_434;
wire n_6_435;
wire n_6_436;
wire n_6_437;
wire n_6_438;
wire n_6_439;
wire n_6_440;
wire n_6_441;
wire n_6_442;
wire n_6_443;
wire n_6_444;
wire n_6_445;
wire n_6_446;
wire n_6_447;
wire n_6_448;
wire n_6_449;
wire n_6_450;
wire n_6_451;
wire n_6_452;
wire n_6_453;
wire n_6_454;
wire n_6_455;
wire n_6_456;
wire n_6_457;
wire n_6_458;
wire n_6_459;
wire n_6_460;
wire n_6_461;
wire n_6_462;
wire n_6_463;
wire n_6_464;
wire n_6_465;
wire n_6_466;
wire n_6_467;
wire n_6_468;
wire n_6_469;
wire n_6_470;
wire n_6_471;
wire n_6_472;
wire n_6_473;
wire n_6_474;
wire n_6_475;
wire n_6_476;
wire n_6_477;
wire n_6_478;
wire n_6_479;
wire n_6_480;
wire n_6_481;
wire n_6_482;
wire n_6_483;
wire n_6_484;
wire n_6_485;
wire n_6_486;
wire n_6_487;
wire n_6_488;
wire n_6_489;
wire n_6_490;
wire n_6_491;
wire n_6_492;
wire n_6_493;
wire n_6_494;
wire n_6_495;
wire n_6_496;
wire n_6_497;
wire n_6_498;
wire n_6_499;
wire n_6_500;
wire n_6_501;
wire n_6_502;
wire n_6_503;
wire n_6_504;
wire n_6_505;
wire n_6_506;
wire n_6_507;
wire n_6_508;
wire n_6_509;
wire n_6_510;
wire n_6_511;
wire n_6_512;
wire n_6_513;
wire n_6_514;
wire n_6_515;
wire n_6_516;
wire n_6_517;
wire n_6_518;
wire n_6_519;
wire n_6_520;
wire n_6_521;
wire n_6_522;
wire n_6_523;
wire n_6_524;
wire n_6_525;
wire n_6_526;
wire n_6_527;
wire n_6_528;
wire n_6_529;
wire n_6_530;
wire n_6_531;
wire n_6_532;
wire n_6_533;
wire n_6_534;
wire n_6_535;
wire n_6_536;
wire n_6_537;
wire n_6_538;
wire n_6_539;
wire n_6_540;
wire n_6_541;
wire n_6_542;
wire n_6_543;
wire n_6_544;
wire n_6_545;
wire n_6_546;
wire n_6_547;
wire n_6_548;
wire n_6_549;
wire n_6_550;
wire n_6_551;
wire n_6_552;
wire n_6_553;
wire n_6_554;
wire n_6_555;
wire n_6_556;
wire n_6_557;
wire n_6_558;
wire n_6_559;
wire n_6_560;
wire n_6_561;
wire n_6_562;
wire n_6_563;
wire n_6_564;
wire n_6_565;
wire n_6_566;
wire n_6_567;
wire n_6_568;
wire n_6_569;
wire n_6_570;
wire n_6_571;
wire n_6_572;
wire n_6_573;
wire n_6_574;
wire n_6_575;
wire n_6_576;
wire n_6_577;
wire n_6_578;
wire n_6_579;
wire n_6_580;
wire n_6_581;
wire n_6_582;
wire n_6_583;
wire n_6_584;
wire n_6_585;
wire n_6_586;
wire n_6_587;
wire n_6_588;
wire n_6_589;
wire n_6_590;
wire n_6_591;
wire n_6_592;
wire n_6_593;
wire n_6_594;
wire n_6_595;
wire n_6_596;
wire n_6_597;
wire n_6_598;
wire n_6_599;
wire n_6_600;
wire n_6_601;
wire n_6_602;
wire n_6_603;
wire n_6_604;
wire n_6_605;
wire n_6_606;
wire n_6_607;
wire n_6_608;
wire n_6_609;
wire n_6_610;
wire n_6_611;
wire n_6_612;
wire n_6_613;
wire n_6_614;
wire n_6_615;
wire n_6_616;
wire n_6_617;
wire n_6_618;
wire n_6_619;
wire n_6_620;
wire n_6_621;
wire n_6_622;
wire n_6_623;
wire n_6_624;
wire n_6_625;
wire n_6_626;
wire n_6_627;
wire n_6_628;
wire n_6_629;
wire n_6_630;
wire n_6_631;
wire n_6_632;
wire n_6_633;
wire n_6_634;
wire n_6_635;
wire n_6_636;
wire n_6_637;
wire n_6_638;
wire n_6_639;
wire n_6_640;
wire n_6_641;
wire n_6_642;
wire n_6_643;
wire n_6_644;
wire n_6_645;
wire n_6_646;
wire n_6_647;
wire n_6_648;
wire n_6_649;
wire n_6_650;
wire n_6_651;
wire n_6_652;
wire n_6_653;
wire n_6_654;
wire n_6_655;
wire n_6_656;
wire n_6_657;
wire n_6_658;
wire n_6_659;
wire n_6_660;
wire n_6_661;
wire n_6_662;
wire n_6_663;
wire n_6_664;
wire n_6_665;
wire n_6_666;
wire n_6_667;
wire n_6_668;
wire n_6_669;
wire n_6_670;
wire n_6_671;
wire n_6_672;
wire n_6_673;
wire n_6_674;
wire n_6_675;
wire n_6_676;
wire n_6_677;
wire n_6_678;
wire n_6_679;
wire n_6_680;
wire n_6_681;
wire n_6_682;
wire n_6_683;
wire n_6_684;
wire n_6_685;
wire n_6_686;
wire n_6_687;
wire n_6_688;
wire n_6_689;
wire n_6_690;
wire n_6_691;
wire n_6_692;
wire n_6_693;
wire n_6_694;
wire n_6_695;
wire n_6_696;
wire n_6_697;
wire n_6_698;
wire n_6_699;
wire n_6_700;
wire n_6_701;
wire n_6_702;
wire n_6_703;
wire n_6_704;
wire n_6_705;
wire n_6_706;
wire n_6_707;
wire n_6_708;
wire n_6_709;
wire n_6_710;
wire n_6_711;
wire n_6_712;
wire n_6_713;
wire n_6_714;
wire n_6_715;
wire n_6_716;
wire n_6_717;
wire n_6_718;
wire n_6_719;
wire n_6_720;
wire n_6_721;
wire n_6_722;
wire n_6_723;
wire n_6_724;
wire n_6_725;
wire n_6_726;
wire n_6_727;
wire n_6_728;
wire n_6_729;
wire n_6_730;
wire n_6_731;
wire n_6_732;
wire n_6_733;
wire n_6_734;
wire n_6_735;
wire n_6_736;
wire n_6_737;
wire n_6_738;
wire n_6_739;
wire n_6_740;
wire n_6_741;
wire n_6_742;
wire n_6_743;
wire n_6_744;
wire n_6_745;
wire n_6_746;
wire n_6_747;
wire n_6_748;
wire n_6_749;
wire n_6_750;
wire n_6_751;
wire n_6_752;
wire n_6_753;
wire n_6_754;
wire n_6_755;
wire n_6_756;
wire n_6_757;
wire n_6_758;
wire n_6_759;
wire n_6_760;
wire n_6_761;
wire n_6_762;
wire n_6_763;
wire n_6_764;
wire n_6_765;
wire n_6_766;
wire n_6_767;
wire n_6_768;
wire n_6_769;
wire n_6_770;
wire n_6_771;
wire n_6_772;
wire n_6_773;
wire n_6_774;
wire n_6_775;
wire n_6_776;
wire n_6_777;
wire n_6_778;
wire n_6_779;
wire n_6_780;
wire n_6_781;
wire n_6_782;
wire n_6_783;
wire n_6_784;
wire n_6_785;
wire n_6_786;
wire n_6_787;
wire n_6_788;
wire n_6_789;
wire n_6_790;
wire n_6_791;
wire n_6_792;
wire n_6_793;
wire n_6_794;
wire n_6_795;
wire n_6_796;
wire n_6_797;
wire n_6_798;
wire n_6_799;
wire n_6_800;
wire n_6_801;
wire n_6_802;
wire n_6_803;
wire n_6_804;
wire n_6_805;
wire n_6_806;
wire n_6_807;
wire n_6_808;
wire n_6_809;
wire n_6_810;
wire n_6_811;
wire n_6_812;
wire n_6_813;
wire n_6_814;
wire n_6_815;
wire n_6_816;
wire n_6_817;
wire n_6_818;
wire n_6_819;
wire n_6_820;
wire n_6_821;
wire n_6_822;
wire n_6_823;
wire n_6_824;
wire n_6_825;
wire n_6_826;
wire n_6_827;
wire n_6_828;
wire n_6_829;
wire n_6_830;
wire n_6_831;
wire n_6_832;
wire n_6_833;
wire n_6_834;
wire n_6_835;
wire n_6_836;
wire n_6_837;
wire n_6_838;
wire n_6_839;
wire n_6_840;
wire n_6_841;
wire n_6_842;
wire n_6_843;
wire n_6_844;
wire n_6_845;
wire n_6_846;
wire n_6_847;
wire n_6_848;
wire n_6_849;
wire n_6_850;
wire n_6_851;
wire n_6_852;
wire n_6_853;
wire n_6_854;
wire n_6_855;
wire n_6_856;
wire n_6_857;
wire n_6_858;
wire n_6_859;
wire n_6_860;
wire n_6_861;
wire n_6_862;
wire n_6_863;
wire n_6_864;
wire n_6_865;
wire n_6_866;
wire n_6_867;
wire n_6_868;
wire n_6_869;
wire n_6_870;
wire n_6_871;
wire n_6_872;
wire n_6_873;
wire n_6_874;
wire n_6_875;
wire n_6_876;
wire n_6_877;
wire n_6_878;
wire n_6_879;
wire n_6_880;
wire n_6_881;
wire n_6_882;
wire n_6_883;
wire n_6_884;
wire n_6_885;
wire n_6_886;
wire n_6_887;
wire n_6_888;
wire n_6_889;
wire n_6_890;
wire n_6_891;
wire n_6_892;
wire n_6_893;
wire n_6_894;
wire n_6_895;
wire n_6_896;
wire n_6_897;
wire n_6_898;
wire n_6_899;
wire n_6_900;
wire n_6_901;
wire n_6_902;
wire n_6_903;
wire n_6_904;
wire n_6_905;
wire n_6_906;
wire n_6_907;
wire n_6_908;
wire n_6_909;
wire n_6_910;
wire n_6_911;
wire n_6_912;
wire n_6_913;
wire n_6_914;
wire n_6_915;
wire n_6_916;
wire n_6_917;
wire n_6_918;
wire n_6_919;
wire n_6_920;
wire n_6_921;
wire n_6_922;
wire n_6_923;
wire n_6_924;
wire n_6_925;
wire n_6_926;
wire n_6_927;
wire n_6_928;
wire n_6_929;
wire n_6_930;
wire n_6_931;
wire n_6_932;
wire n_6_933;
wire n_6_934;
wire n_6_935;
wire n_6_936;
wire n_6_937;
wire n_6_938;
wire n_6_939;
wire n_6_940;
wire n_6_941;
wire n_6_942;
wire n_6_943;
wire n_6_944;
wire n_6_945;
wire n_6_946;
wire n_6_947;
wire n_6_948;
wire n_6_949;
wire n_6_950;
wire n_6_951;
wire n_6_952;
wire n_6_953;
wire n_6_954;
wire n_6_955;
wire n_6_956;
wire n_6_957;
wire n_6_958;
wire n_6_959;
wire n_6_960;
wire n_6_961;
wire n_6_962;
wire n_6_963;
wire n_6_964;
wire n_6_965;
wire n_6_966;
wire n_6_967;
wire n_6_968;
wire n_6_969;
wire n_6_970;
wire n_6_971;
wire n_6_972;
wire n_6_973;
wire n_6_974;
wire n_6_975;
wire n_6_976;
wire n_6_977;
wire n_6_978;
wire n_6_979;
wire n_6_980;
wire n_6_981;
wire n_6_982;
wire n_6_983;
wire n_6_984;
wire n_6_985;
wire n_6_986;
wire n_6_987;
wire n_6_988;
wire n_6_989;
wire n_6_990;
wire n_6_991;
wire n_6_992;
wire n_6_993;
wire n_6_994;
wire n_6_995;
wire n_6_996;
wire n_6_997;
wire n_6_998;
wire n_6_999;
wire n_6_1000;
wire n_6_1001;
wire n_6_1002;
wire n_6_1003;
wire n_6_1004;
wire n_6_1005;
wire n_6_1006;
wire n_6_1007;
wire n_6_1008;
wire n_6_1009;
wire n_6_1010;
wire n_6_1011;
wire n_6_1012;
wire n_6_1013;
wire n_6_1014;
wire n_6_1015;
wire n_6_1016;
wire n_6_1017;
wire n_6_1018;
wire n_6_1019;
wire n_6_1020;
wire n_6_1021;
wire n_6_1022;
wire n_6_1023;
wire n_6_1024;
wire n_6_1025;
wire n_6_1026;
wire n_6_1027;
wire n_6_1028;
wire n_6_1029;
wire n_6_1030;
wire n_6_1031;
wire n_6_1032;
wire n_6_1033;
wire n_6_1034;
wire n_6_1035;
wire n_6_1036;
wire n_6_1037;
wire n_6_1038;
wire n_6_1039;
wire n_6_1040;
wire n_6_1041;
wire n_6_1042;
wire n_6_1043;
wire n_6_1044;
wire n_6_1045;
wire n_6_1046;
wire n_6_1047;
wire n_6_1048;
wire n_6_1049;
wire n_6_1050;
wire n_6_1051;
wire n_6_1052;
wire n_6_1053;
wire n_6_1054;
wire n_6_1055;
wire n_6_1056;
wire n_6_1057;
wire n_6_1058;
wire n_6_1059;
wire n_6_1060;
wire n_6_1061;
wire n_6_1062;
wire n_6_1063;
wire n_6_1064;
wire n_6_1065;
wire n_6_1066;
wire n_6_1067;
wire n_6_1068;
wire n_6_1069;
wire n_6_1070;
wire n_6_1071;
wire n_6_1072;
wire n_6_1073;
wire n_6_1074;
wire n_6_1075;
wire n_6_1076;
wire n_6_1077;
wire n_6_1078;
wire n_6_1079;
wire n_6_1080;
wire n_6_1081;
wire n_6_1082;
wire n_6_1083;
wire n_6_1084;
wire n_6_1085;
wire n_6_1086;
wire n_6_1087;
wire n_6_1088;
wire n_6_1089;
wire n_6_1090;
wire n_6_1091;
wire n_6_1092;
wire n_6_1093;
wire n_6_1094;
wire n_6_1095;
wire n_6_1096;
wire n_6_1097;
wire n_6_1098;
wire n_6_1099;
wire n_6_1100;
wire n_6_1101;
wire n_6_1102;
wire n_6_1103;
wire n_6_1104;
wire n_6_1105;
wire n_6_1106;
wire n_6_1107;
wire n_6_1108;
wire n_6_1109;
wire n_6_1110;
wire n_6_1111;
wire n_6_1112;
wire n_6_1113;
wire n_6_1114;
wire n_6_1115;
wire n_6_1116;
wire n_6_1117;
wire n_6_1118;
wire n_6_1119;
wire n_6_1120;
wire n_6_1121;
wire n_6_1122;
wire n_6_1123;
wire n_6_1124;
wire n_6_1125;
wire n_6_1126;
wire n_6_1127;
wire n_6_1128;
wire n_6_1129;
wire n_6_1130;
wire n_6_1131;
wire n_6_1132;
wire n_6_1133;
wire n_6_1134;
wire n_6_1135;
wire n_6_1136;
wire n_6_1137;
wire n_6_1138;
wire n_6_1139;
wire n_6_1140;
wire n_6_1141;
wire n_6_1142;
wire n_6_1143;
wire n_6_1144;
wire n_6_1145;
wire n_6_1146;
wire n_6_1147;
wire n_6_1148;
wire n_6_1149;
wire n_6_1150;
wire n_6_1151;
wire n_6_1152;
wire n_6_1153;
wire n_6_1154;
wire n_6_1155;
wire n_6_1156;
wire n_6_1157;
wire n_6_1158;
wire n_6_1159;
wire n_6_1160;
wire n_6_1161;
wire n_6_1162;
wire n_6_1163;
wire n_6_1164;
wire n_6_1165;
wire n_6_1166;
wire n_6_1167;
wire n_6_1168;
wire n_6_1169;
wire n_6_1170;
wire n_6_1171;
wire n_6_1172;
wire n_6_1173;
wire n_6_1174;
wire n_6_1175;
wire n_6_1176;
wire n_6_1177;
wire n_6_1178;
wire n_6_1179;
wire n_6_1180;
wire n_6_1181;
wire n_6_1182;
wire n_6_1183;
wire n_6_1184;
wire n_6_1185;
wire n_6_1186;
wire n_6_1187;
wire n_6_1188;
wire n_6_1189;
wire n_6_1190;
wire n_6_1191;
wire n_6_1192;
wire n_6_1193;
wire n_6_1194;
wire n_6_1195;
wire n_6_1196;
wire n_6_1197;
wire n_6_1198;
wire n_6_1199;
wire n_6_1200;
wire n_6_1201;
wire n_6_1202;
wire n_6_1203;
wire n_6_1204;
wire n_6_1205;
wire n_6_1206;
wire n_6_1207;
wire n_6_1208;
wire n_6_1209;
wire n_6_1210;
wire n_6_1211;
wire n_6_1212;
wire n_6_1213;
wire n_6_1214;
wire n_6_1215;
wire n_6_1216;
wire n_6_1217;
wire n_6_1218;
wire n_6_1219;
wire n_6_1220;
wire n_6_1221;
wire n_6_1222;
wire n_6_1223;
wire n_6_1224;
wire n_6_1225;
wire n_6_1226;
wire n_6_1227;
wire n_6_1228;
wire n_6_1229;
wire n_6_1230;
wire n_6_1231;
wire n_6_1232;
wire n_6_1233;
wire n_6_1234;
wire n_6_1235;
wire n_6_1236;
wire n_6_1237;
wire n_6_1238;
wire n_6_1239;
wire n_6_1240;
wire n_6_1241;
wire n_6_1242;
wire n_6_1243;
wire n_6_1244;
wire n_6_1245;
wire n_6_1246;
wire n_6_1247;
wire n_6_1248;
wire n_6_1249;
wire n_6_1250;
wire n_6_1251;
wire n_6_1252;
wire n_6_1253;
wire n_6_1254;
wire n_6_1255;
wire n_6_1256;
wire n_6_1257;
wire n_6_1258;
wire n_6_1259;
wire n_6_1260;
wire n_6_1261;
wire n_6_1262;
wire n_6_1263;
wire n_6_1264;
wire n_6_1265;
wire n_6_1266;
wire n_6_1267;
wire n_6_1268;
wire n_6_1269;
wire n_6_1270;
wire n_6_1271;
wire n_6_1272;
wire n_6_1273;
wire n_6_1274;
wire n_6_1275;
wire n_6_1276;
wire n_6_1277;
wire n_6_1278;
wire n_6_1279;
wire n_6_1280;
wire n_6_1281;
wire n_6_1282;
wire n_6_1283;
wire n_6_1284;
wire n_6_1285;
wire n_6_1286;
wire n_6_1287;
wire n_6_1288;
wire n_6_1289;
wire n_6_1290;
wire n_6_1291;
wire n_6_1292;
wire n_6_1293;
wire n_6_1294;
wire n_6_1295;
wire n_6_1296;
wire n_6_1297;
wire n_6_1298;
wire n_6_1299;
wire n_6_1300;
wire n_6_1301;
wire n_6_1302;
wire n_6_1303;
wire n_6_1304;
wire n_6_1305;
wire n_6_1306;
wire n_6_1307;
wire n_6_1308;
wire n_6_1309;
wire n_6_1310;
wire n_6_1311;
wire n_6_1312;
wire n_6_1313;
wire n_6_1314;
wire n_6_1315;
wire n_6_1316;
wire n_6_1317;
wire n_6_1318;
wire n_6_1319;
wire n_6_1320;
wire n_6_1321;
wire n_6_1322;
wire n_6_1323;
wire n_6_1324;
wire n_6_1325;
wire n_6_1326;
wire n_6_1327;
wire n_6_1328;
wire n_6_1329;
wire n_6_1330;
wire n_6_1331;
wire n_6_1332;
wire n_6_1333;
wire n_6_1334;
wire n_6_1335;
wire n_6_1336;
wire n_6_1337;
wire n_6_1338;
wire n_6_1339;
wire n_6_1340;
wire n_6_1341;
wire n_6_1342;
wire n_6_1343;
wire n_6_1344;
wire n_6_1345;
wire n_6_1346;
wire n_6_1347;
wire n_6_1348;
wire n_6_1349;
wire n_6_1350;
wire n_6_1351;
wire n_6_1352;
wire n_6_1353;
wire n_6_1354;
wire n_6_1355;
wire n_6_1356;
wire n_6_1357;
wire n_6_1358;
wire n_6_1359;
wire n_6_1360;
wire n_6_1361;
wire n_6_1362;
wire n_6_1363;
wire n_6_1364;
wire n_6_1365;
wire n_6_1366;
wire n_6_1367;
wire n_6_1368;
wire n_6_1369;
wire n_6_1370;
wire n_6_1371;
wire n_6_1372;
wire n_6_1373;
wire n_6_1374;
wire n_6_1375;
wire n_6_1376;
wire n_6_1377;
wire n_6_1378;
wire n_6_1379;
wire n_6_1380;
wire n_6_1381;
wire n_6_1382;
wire n_6_1383;
wire n_6_1384;
wire n_6_1385;
wire n_6_1386;
wire n_6_1387;
wire n_6_1388;
wire n_6_1389;
wire n_6_1390;
wire n_6_1391;
wire n_6_1392;
wire n_6_1393;
wire n_6_1394;
wire n_6_1395;
wire n_6_1396;
wire n_6_1397;
wire n_6_1398;
wire n_6_1399;
wire n_6_1400;
wire n_6_1401;
wire n_6_1402;
wire n_6_1403;
wire n_6_1404;
wire n_6_1405;
wire n_6_1406;
wire n_6_1407;
wire n_6_1408;
wire n_6_1409;
wire n_6_1410;
wire n_6_1411;
wire n_6_1412;
wire n_6_1413;
wire n_6_1414;
wire n_6_1415;
wire n_6_1416;
wire n_6_1417;
wire n_6_1418;
wire n_6_1419;
wire n_6_1420;
wire n_6_1421;
wire n_6_1422;
wire n_6_1423;
wire n_6_1424;
wire n_6_1425;
wire n_6_1426;
wire n_6_1427;
wire n_6_1428;
wire n_6_1429;
wire n_6_1430;
wire n_6_1431;
wire n_6_1432;
wire n_6_1433;
wire n_6_1434;
wire n_6_1435;
wire n_6_1436;
wire n_6_1437;
wire n_6_1438;
wire n_6_1439;
wire n_6_1440;
wire n_6_1441;
wire n_6_1442;
wire n_6_1443;
wire n_6_1444;
wire n_6_1445;
wire n_6_1446;
wire n_6_1447;
wire n_6_1448;
wire n_6_1449;
wire n_6_1450;
wire n_6_1451;
wire n_6_1452;
wire n_6_1453;
wire n_6_1454;
wire n_6_1455;
wire n_6_1456;
wire n_6_1457;
wire n_6_1458;
wire n_6_1459;
wire n_6_1460;
wire n_6_1461;
wire n_6_1462;
wire n_6_1463;
wire n_6_1464;
wire n_6_1465;
wire n_6_1466;
wire n_6_1467;
wire n_6_1468;
wire n_6_1469;
wire n_6_1470;
wire n_6_1471;
wire n_6_1472;
wire n_6_1473;
wire n_6_1474;
wire n_6_1475;
wire n_6_1476;
wire n_6_1477;
wire n_6_1478;
wire n_6_1479;
wire n_6_1480;
wire n_6_1481;
wire n_6_1482;
wire n_6_1483;
wire n_6_1484;
wire n_6_1485;
wire n_6_1486;
wire n_6_1487;
wire n_6_1488;
wire n_6_1489;
wire n_6_1490;
wire n_6_1491;
wire n_6_1492;
wire n_6_1493;
wire n_6_1494;
wire n_6_1495;
wire n_6_1496;
wire n_6_1497;
wire n_6_1498;
wire n_6_1499;
wire n_6_1500;
wire n_6_1501;
wire n_6_1502;
wire n_6_1503;
wire n_6_1504;
wire n_6_1505;
wire n_6_1506;
wire n_6_1507;
wire n_6_1508;
wire n_6_1509;
wire n_6_1510;
wire n_6_1511;
wire n_6_1512;
wire n_6_1513;
wire n_6_1514;
wire n_6_1515;
wire n_6_1516;
wire n_6_1517;
wire n_6_1518;
wire n_6_1519;
wire n_6_1520;
wire n_6_1521;
wire n_6_1522;
wire n_6_1523;
wire n_6_1524;
wire n_6_1525;
wire n_6_1526;
wire n_6_1527;
wire n_6_1528;
wire n_6_1529;
wire n_6_1530;
wire n_6_1531;
wire n_6_1532;
wire n_6_1533;
wire n_6_1534;
wire n_6_1535;
wire n_6_1536;
wire n_6_1537;
wire n_6_1538;
wire n_6_1539;
wire n_6_1540;
wire n_6_1541;
wire n_6_1542;
wire n_6_1543;
wire n_6_1544;
wire n_6_1545;
wire n_6_1546;
wire n_6_1547;
wire n_6_1548;
wire n_6_1549;
wire n_6_1550;
wire n_6_1551;
wire n_6_1552;
wire n_6_1553;
wire n_6_1554;
wire n_6_1555;
wire n_6_1556;
wire n_6_1557;
wire n_6_1558;
wire n_6_1559;
wire n_6_1560;
wire n_6_1561;
wire n_6_1562;
wire n_6_1563;
wire n_6_1564;
wire n_6_1565;
wire n_6_1566;
wire n_6_1567;
wire n_6_1568;
wire n_6_1569;
wire n_6_1570;
wire n_6_1571;
wire n_6_1572;
wire n_6_1573;
wire n_6_1574;
wire n_6_1575;
wire n_6_1576;
wire n_6_1577;
wire n_6_1578;
wire n_6_1579;
wire n_6_1580;
wire n_6_1581;
wire n_6_1582;
wire n_6_1583;
wire n_6_1584;
wire n_6_1585;
wire n_6_1586;
wire n_6_1587;
wire n_6_1588;
wire n_6_1589;
wire n_6_1590;
wire n_6_1591;
wire n_6_1592;
wire n_6_1593;
wire n_6_1594;
wire n_6_1595;
wire n_6_1596;
wire n_6_1597;
wire n_6_1598;
wire n_6_1599;
wire n_6_1600;
wire n_6_1601;
wire n_6_1602;
wire n_6_1603;
wire n_6_1604;
wire n_6_1605;
wire n_6_1606;
wire n_6_1607;
wire n_6_1608;
wire n_6_1609;
wire n_6_1610;
wire n_6_1611;
wire n_6_1612;
wire n_6_1613;
wire n_6_1614;
wire n_6_1615;
wire n_6_1616;
wire n_6_1617;
wire n_6_1618;
wire n_6_1619;
wire n_6_1620;
wire n_6_1621;
wire n_6_1622;
wire n_6_1623;
wire n_6_1624;
wire n_6_1625;
wire n_6_1626;
wire n_6_1627;
wire n_6_1628;
wire n_6_1629;
wire n_6_1630;
wire n_6_1631;
wire n_6_1632;
wire n_6_1633;
wire n_6_1634;
wire n_6_1635;
wire n_6_1636;
wire n_6_1637;
wire n_6_1638;
wire n_6_1639;
wire n_6_1640;
wire n_6_1641;
wire n_6_1642;
wire n_6_1643;
wire n_6_1644;
wire n_6_1645;
wire n_6_1646;
wire n_6_1647;
wire n_6_1648;
wire n_6_1649;
wire n_6_1650;
wire n_6_1651;
wire n_6_1652;
wire n_6_1653;
wire n_6_1654;
wire n_6_1655;
wire n_6_1656;
wire n_6_1657;
wire n_6_1658;
wire n_6_1659;
wire n_6_1660;
wire n_6_1661;
wire n_6_1662;
wire n_6_1663;
wire n_6_1664;
wire n_6_1665;
wire n_6_1666;
wire n_6_1667;
wire n_6_1668;
wire n_6_1669;
wire n_6_1670;
wire n_6_1671;
wire n_6_1672;
wire n_6_1673;
wire n_6_1674;
wire n_6_1675;
wire n_6_1676;
wire n_6_1677;
wire n_6_1678;
wire n_6_1679;
wire n_6_1680;
wire n_6_1681;
wire n_6_1682;
wire n_6_1683;
wire n_6_1684;
wire n_6_1685;
wire n_6_1686;
wire n_6_1687;
wire n_6_1688;
wire n_6_1689;
wire n_6_1690;
wire n_6_1691;
wire n_6_1692;
wire n_6_1693;
wire n_6_1694;
wire n_6_1695;
wire n_6_1696;
wire n_6_1697;
wire n_6_1698;
wire n_6_1699;
wire n_6_1700;
wire n_6_1701;
wire n_6_1702;
wire n_6_1703;
wire n_6_1704;
wire n_6_1705;
wire n_6_1706;
wire n_6_1707;
wire n_6_1708;
wire n_6_1709;
wire n_6_1710;
wire n_6_1711;
wire n_6_1712;
wire n_6_1713;
wire n_6_1714;
wire n_6_1715;
wire n_6_1716;
wire n_6_1717;
wire n_6_1718;
wire n_6_1719;
wire n_6_1720;
wire n_6_1721;
wire n_6_1722;
wire n_6_1723;
wire n_6_1724;
wire n_6_1725;
wire n_6_1726;
wire n_6_1727;
wire n_6_1728;
wire n_6_1729;
wire n_6_1730;
wire n_6_1731;
wire n_6_1732;
wire n_6_1733;
wire n_6_1734;
wire n_6_1735;
wire n_6_1736;
wire n_6_1737;
wire n_6_1738;
wire n_6_1739;
wire n_6_1740;
wire n_6_1741;
wire n_6_1742;
wire n_6_1743;
wire n_6_1744;
wire n_6_1745;
wire n_6_1746;
wire n_6_1747;
wire n_6_1748;
wire n_6_1749;
wire n_6_1750;
wire n_6_1751;
wire n_6_1752;
wire n_6_1753;
wire n_6_1754;
wire n_6_1755;
wire n_6_1756;
wire n_6_1757;
wire n_6_1758;
wire n_6_1759;
wire n_6_1760;
wire n_6_1761;
wire n_6_1762;
wire n_6_1763;
wire n_6_1764;
wire n_6_1765;
wire n_6_1766;
wire n_6_1767;
wire n_6_1768;
wire n_6_1769;
wire n_6_1770;
wire n_6_1771;
wire n_6_1772;
wire n_6_1773;
wire n_6_1774;
wire n_6_1775;
wire n_6_1776;
wire n_6_1777;
wire n_6_1778;
wire n_6_1779;
wire n_6_1780;
wire n_6_1781;
wire n_6_1782;
wire n_6_1783;
wire n_6_1784;
wire n_6_1785;
wire n_6_1786;
wire n_6_1787;
wire n_6_1788;
wire n_6_1789;
wire n_6_1790;
wire n_6_1791;
wire n_6_1792;
wire n_6_1793;
wire n_6_1794;
wire n_6_1795;
wire n_6_1796;
wire n_6_1797;
wire n_6_1798;
wire n_6_1799;
wire n_6_1800;
wire n_6_1801;
wire n_6_1802;
wire n_6_1803;
wire n_6_1804;
wire n_6_1805;
wire n_6_1806;
wire n_6_1807;
wire n_6_1808;
wire n_6_1809;
wire n_6_1810;
wire n_6_1811;
wire n_6_1812;
wire n_6_1813;
wire n_6_1814;
wire n_6_1815;
wire n_6_1816;
wire n_6_1817;
wire n_6_1818;
wire n_6_1819;
wire n_6_1820;
wire n_6_1821;
wire n_6_1822;
wire n_6_1823;
wire n_6_1824;
wire n_6_1825;
wire n_6_1826;
wire n_6_1827;
wire n_6_1828;
wire n_6_1829;
wire n_6_1830;
wire n_6_1831;
wire n_6_1832;
wire n_6_1833;
wire n_6_1834;
wire n_6_1835;
wire n_6_1836;
wire n_6_1837;
wire n_6_1838;
wire n_6_1839;
wire n_6_1840;
wire n_6_1841;
wire n_6_1842;
wire n_6_1843;
wire n_6_1844;
wire n_6_1845;
wire n_6_1846;
wire n_6_1847;
wire n_6_1848;
wire n_6_1849;
wire n_6_1850;
wire n_6_1851;
wire n_6_1852;
wire n_6_1853;
wire n_6_1854;
wire n_6_1855;
wire n_6_1856;
wire n_6_1857;
wire n_6_1858;
wire n_6_1859;
wire n_6_1860;
wire n_6_1861;
wire n_6_1862;
wire n_6_1863;
wire n_6_1864;
wire n_6_1865;
wire n_6_1866;
wire n_6_1867;
wire n_6_1868;
wire n_6_1869;
wire n_6_1870;
wire n_6_1871;
wire n_6_1872;
wire n_6_1873;
wire n_6_1874;
wire n_6_1875;
wire n_6_1876;
wire n_6_1877;
wire n_6_1878;
wire n_6_1879;
wire n_6_1880;
wire n_6_1881;
wire n_6_1882;
wire n_6_1883;
wire n_6_1884;
wire n_6_1885;
wire n_6_1886;
wire n_6_1887;
wire n_6_1888;
wire n_6_1889;
wire n_6_1890;
wire n_6_1891;
wire n_6_1892;
wire n_6_1893;
wire n_6_1894;
wire n_6_1895;
wire n_6_1896;
wire n_6_1897;
wire n_6_1898;
wire n_6_1899;
wire n_6_1900;
wire n_6_1901;
wire n_6_1902;
wire n_6_1903;
wire n_6_1904;
wire n_6_1905;
wire n_6_1906;
wire n_6_1907;
wire n_6_1908;
wire n_6_1909;
wire n_6_1910;
wire n_6_1911;
wire n_6_1912;
wire n_6_1913;
wire n_6_1914;
wire n_6_1915;
wire n_6_1916;
wire n_6_1917;
wire n_6_1918;
wire n_6_1919;
wire n_6_1920;
wire n_6_1921;
wire n_6_1922;
wire n_6_1923;
wire n_6_1924;
wire n_6_1925;
wire n_6_1926;
wire n_6_1927;
wire n_6_1928;
wire n_6_1929;
wire n_6_1930;
wire n_6_1931;
wire n_6_1932;
wire n_6_1933;
wire n_6_1934;
wire n_6_1935;
wire n_6_1936;
wire n_6_1937;
wire n_6_1938;
wire n_6_1939;
wire n_6_1940;
wire n_6_1941;
wire n_6_1942;
wire n_6_1943;
wire n_6_1944;
wire n_6_1945;
wire n_6_1946;
wire n_6_1947;
wire n_6_1948;
wire n_6_1949;
wire n_6_1950;
wire n_6_1951;
wire n_6_1952;
wire n_6_1953;
wire n_6_1954;
wire n_6_1955;
wire n_6_1956;
wire n_6_1957;
wire n_6_1958;
wire n_6_1959;
wire n_6_1960;
wire n_6_1961;
wire n_6_1962;
wire n_6_1963;
wire n_6_1964;
wire n_6_1965;
wire n_6_1966;
wire n_6_1967;
wire n_6_1968;
wire n_6_1969;
wire n_6_1970;
wire n_6_1971;
wire n_6_1972;
wire n_6_1973;
wire n_6_1974;
wire n_6_1975;
wire n_6_1976;
wire n_6_1977;
wire n_6_1978;
wire n_6_1979;
wire n_6_1980;
wire n_6_1981;
wire n_6_1982;
wire n_6_1_0;
wire n_6_1_1;
wire n_6_1_2;
wire n_6_1_3;
wire n_6_1_4;
wire n_6_1_5;
wire n_6_1_6;
wire n_6_1_7;
wire n_6_1_8;
wire n_6_1_9;
wire n_6_1_10;
wire n_6_1_11;
wire n_6_1_12;
wire n_6_1_13;
wire n_6_1_14;
wire n_6_1_15;
wire n_6_1_16;
wire n_6_1_17;
wire n_6_1_18;
wire n_6_1_19;
wire n_6_1_20;
wire n_6_1_21;
wire n_6_1_22;
wire n_6_1_23;
wire n_6_1_24;
wire n_6_1_25;
wire n_6_1_26;
wire n_6_1_27;
wire n_6_1_28;
wire n_6_1_29;
wire n_6_1_30;
wire n_6_1_31;
wire n_6_1_32;
wire n_6_1_33;
wire n_6_1_34;
wire n_6_1_35;
wire n_6_1_36;
wire n_6_1_37;
wire n_6_1_38;
wire n_6_1_39;
wire n_6_1_40;
wire n_6_1_41;
wire n_6_1_42;
wire n_6_1_43;
wire n_6_1_44;
wire n_6_1_45;
wire n_6_1_46;
wire n_6_1_47;
wire n_6_1_48;
wire n_6_1_49;
wire n_6_1_50;
wire n_6_1_51;
wire n_6_1_52;
wire n_6_1_53;
wire n_6_1_54;
wire n_6_1_55;
wire slo__sro_n13037;
wire slo___n13086;
wire n_6_1_58;
wire slo__sro_n33596;
wire slo__mro_n33300;
wire sgo__sro_n1602;
wire n_6_1_62;
wire n_6_1_63;
wire n_6_1_64;
wire n_6_1_65;
wire n_6_1983;
wire n_6_1_66;
wire n_6_1984;
wire n_6_1_67;
wire n_6_1985;
wire n_6_1_68;
wire n_6_1986;
wire n_6_1_69;
wire n_6_1987;
wire n_6_1_70;
wire n_6_1988;
wire slo__sro_n6479;
wire n_6_1989;
wire slo__sro_n11595;
wire n_6_1990;
wire n_6_1_73;
wire CLOCK_slo__sro_n60603;
wire n_6_1_74;
wire n_6_1992;
wire slo__sro_n36835;
wire n_6_1993;
wire CLOCK_slo__n57293;
wire n_6_1994;
wire n_6_1_77;
wire n_6_1995;
wire n_6_1_78;
wire n_6_1996;
wire n_6_1_79;
wire n_6_1997;
wire CLOCK_slo__sro_n51852;
wire n_6_1998;
wire n_6_1_81;
wire n_6_1999;
wire n_6_1_82;
wire n_6_2000;
wire n_6_1_83;
wire n_6_2001;
wire n_6_1_84;
wire n_6_2002;
wire n_6_1_85;
wire n_6_2003;
wire n_6_1_86;
wire n_6_2004;
wire n_6_1_87;
wire n_6_1_88;
wire n_6_2006;
wire slo__n39284;
wire n_6_2007;
wire n_6_1_90;
wire slo__sro_n27582;
wire n_6_2009;
wire slo__sro_n27391;
wire n_6_2010;
wire n_6_1_93;
wire n_6_2011;
wire n_6_1_94;
wire n_6_2012;
wire n_6_1_95;
wire n_6_2013;
wire n_6_1_96;
wire n_6_1_97;
wire n_6_1_98;
wire n_6_1_99;
wire n_6_1_100;
wire n_6_2014;
wire n_6_1_101;
wire n_6_2015;
wire n_6_1_102;
wire n_6_2016;
wire n_6_1_103;
wire n_6_2017;
wire slo__sro_n29067;
wire n_6_2018;
wire slo__sro_n29362;
wire n_6_2019;
wire CLOCK_slo__sro_n61961;
wire slo__sro_n28774;
wire n_6_1_107;
wire n_6_2021;
wire CLOCK_slo__sro_n54487;
wire n_6_2022;
wire n_6_1_109;
wire n_6_2023;
wire slo__sro_n10712;
wire n_6_2024;
wire slo__sro_n10380;
wire n_6_2025;
wire n_6_1_112;
wire n_6_2026;
wire slo__sro_n6480;
wire n_6_2027;
wire slo__sro_n6828;
wire CLOCK_sgo__sro_n47136;
wire n_6_1_115;
wire CLOCK_slo__sro_n62531;
wire slo__sro_n15554;
wire spw__n68416;
wire n_6_1_117;
wire n_6_2031;
wire n_6_1_118;
wire n_6_2032;
wire CLOCK_slo__sro_n55687;
wire n_6_2033;
wire n_6_1_120;
wire n_6_2034;
wire n_6_1_121;
wire n_6_2035;
wire slo__sro_n13354;
wire n_6_2036;
wire n_6_1_123;
wire n_6_2037;
wire n_6_1_124;
wire n_6_1_125;
wire n_6_2039;
wire slo__sro_n10838;
wire n_6_2040;
wire n_6_1_127;
wire n_6_2041;
wire slo__sro_n22623;
wire n_6_2042;
wire n_6_1_129;
wire n_6_2043;
wire n_6_1_130;
wire n_6_2044;
wire n_6_1_131;
wire n_6_1_132;
wire n_6_1_133;
wire n_6_1_134;
wire n_6_1_135;
wire n_6_2045;
wire n_6_1_136;
wire n_6_2046;
wire n_6_1_137;
wire n_6_2047;
wire n_6_1_138;
wire n_6_2048;
wire n_6_1_139;
wire n_6_2049;
wire slo__n39452;
wire n_6_2050;
wire n_6_1_141;
wire n_6_2051;
wire slo__sro_n39795;
wire n_6_2052;
wire n_6_1_143;
wire n_6_2053;
wire slo__sro_n4672;
wire n_6_2054;
wire n_6_1_145;
wire n_6_2055;
wire n_6_1_146;
wire n_6_2056;
wire slo__sro_n15670;
wire n_6_2057;
wire n_6_1_148;
wire n_6_2058;
wire slo__sro_n15657;
wire CLOCK_slo__sro_n48959;
wire n_6_1_150;
wire n_6_2060;
wire slo__sro_n13019;
wire n_6_2061;
wire slo__n14771;
wire n_6_2062;
wire slo__n13290;
wire slo__n39406;
wire n_6_1_154;
wire n_6_2064;
wire n_6_1_155;
wire n_6_2065;
wire slo__sro_n35272;
wire n_6_2066;
wire CLOCK_slo__sro_n57156;
wire n_6_2067;
wire n_6_1_158;
wire n_6_2068;
wire slo__sro_n13370;
wire n_6_2069;
wire n_6_1_160;
wire n_6_2070;
wire CLOCK_slo__sro_n52669;
wire n_6_2071;
wire n_6_1_162;
wire n_6_2072;
wire n_6_1_163;
wire n_6_2073;
wire n_6_1_164;
wire n_6_2074;
wire n_6_1_165;
wire n_6_2075;
wire n_6_1_166;
wire n_6_1_167;
wire n_6_1_168;
wire n_6_1_169;
wire n_6_1_170;
wire n_6_2076;
wire n_6_1_171;
wire n_6_2077;
wire n_6_1_172;
wire n_6_2078;
wire slo__sro_n30285;
wire n_6_2079;
wire slo__sro_n6653;
wire n_6_2080;
wire slo__sro_n9534;
wire n_6_2081;
wire slo__sro_n10769;
wire n_6_2082;
wire CLOCK_slo__sro_n54489;
wire n_6_2083;
wire CLOCK_slo__sro_n54567;
wire CLOCK_slo__sro_n51260;
wire slo__sro_n31052;
wire n_6_2085;
wire n_6_1_180;
wire n_6_2086;
wire slo__n14486;
wire n_6_2087;
wire n_6_1_182;
wire n_6_2088;
wire slo__sro_n5963;
wire n_6_2089;
wire slo__n36492;
wire n_6_2090;
wire slo__n13394;
wire slo__sro_n37453;
wire slo__sro_n14274;
wire n_6_2092;
wire n_6_1_187;
wire n_6_2093;
wire slo__sro_n11578;
wire n_6_2094;
wire slo__sro_n14590;
wire n_6_2095;
wire slo__sro_n20612;
wire drc_ipo_n26607;
wire n_6_1_191;
wire n_6_2097;
wire slo__sro_n11746;
wire n_6_2098;
wire slo__sro_n14179;
wire n_6_2099;
wire slo__sro_n30017;
wire n_6_2100;
wire slo__sro_n33814;
wire n_6_2101;
wire n_6_1_196;
wire n_6_2102;
wire slo__sro_n20259;
wire n_6_2103;
wire slo__sro_n13262;
wire n_6_1_199;
wire n_6_2105;
wire n_6_1_200;
wire n_6_2106;
wire n_6_1_201;
wire n_6_1_202;
wire n_6_1_203;
wire n_6_1_204;
wire n_6_1_205;
wire n_6_2107;
wire n_6_1_206;
wire n_6_2108;
wire n_6_1_207;
wire n_6_2109;
wire n_6_1_208;
wire n_6_2110;
wire slo__sro_n31670;
wire n_6_2111;
wire n_6_1_210;
wire n_6_2112;
wire CLOCK_slo__sro_n51619;
wire n_6_2113;
wire n_6_1_212;
wire n_6_2114;
wire n_6_1_213;
wire n_6_2115;
wire slo__sro_n10770;
wire n_6_2116;
wire slo__sro_n5907;
wire n_6_2117;
wire slo__sro_n15586;
wire slo__mro_n33015;
wire n_6_1_217;
wire n_6_2119;
wire n_6_1_218;
wire n_6_2120;
wire CLOCK_slo__sro_n49853;
wire n_6_2121;
wire slo__n18465;
wire n_6_2122;
wire n_6_1_221;
wire n_6_2123;
wire n_6_1_222;
wire n_6_2124;
wire n_6_1_223;
wire n_6_2125;
wire n_6_1_224;
wire n_6_2126;
wire slo__n15402;
wire n_6_2127;
wire n_6_1_226;
wire n_6_2128;
wire slo__sro_n4880;
wire CLOCK_sgo__sro_n47824;
wire slo__sro_n6519;
wire n_6_2130;
wire slo__sro_n22325;
wire CLOCK_slo__n54206;
wire n_6_2132;
wire n_6_1_231;
wire n_6_2133;
wire slo__sro_n35163;
wire n_6_2134;
wire n_6_1_233;
wire n_6_2135;
wire slo__sro_n32202;
wire n_6_2136;
wire n_6_1_235;
wire n_6_2137;
wire n_6_1_236;
wire n_6_1_237;
wire n_6_1_238;
wire n_6_1_239;
wire n_6_1_240;
wire n_6_2138;
wire n_6_1_241;
wire n_6_2139;
wire n_6_1_242;
wire n_6_2140;
wire n_6_1_243;
wire n_6_2141;
wire n_6_1_244;
wire n_6_2142;
wire n_6_1_245;
wire n_6_2143;
wire slo__sro_n18403;
wire n_6_2144;
wire slo__sro_n32485;
wire n_6_2145;
wire n_6_1_248;
wire n_6_2146;
wire slo__sro_n19079;
wire n_6_2147;
wire slo__sro_n15830;
wire n_6_2148;
wire slo__sro_n12556;
wire n_6_2149;
wire n_6_1_252;
wire slo__n38218;
wire n_6_2151;
wire CLOCK_spw__n65836;
wire n_6_2152;
wire slo___n13100;
wire n_6_2153;
wire slo__sro_n3748;
wire n_6_2154;
wire n_6_1_257;
wire n_6_2155;
wire CLOCK_sgo__sro_n47663;
wire opt_ipo_n26244;
wire n_6_1_259;
wire n_6_2157;
wire n_6_1_260;
wire n_6_2158;
wire slo__sro_n7037;
wire n_6_2159;
wire CLOCK_slo__n50780;
wire n_6_2160;
wire slo__sro_n33755;
wire n_6_2161;
wire slo__sro_n15700;
wire n_6_2162;
wire slo__sro_n15684;
wire n_6_2163;
wire slo__sro_n34621;
wire n_6_2164;
wire n_6_1_267;
wire n_6_2165;
wire n_6_1_268;
wire n_6_2166;
wire slo__sro_n27837;
wire n_6_2167;
wire n_6_1_270;
wire n_6_2168;
wire CLOCK_slo__sro_n58341;
wire n_6_1_272;
wire n_6_1_273;
wire n_6_1_274;
wire n_6_1_275;
wire n_6_2169;
wire n_6_1_276;
wire n_6_2170;
wire slo__n36345;
wire n_6_2171;
wire slo__sro_n20509;
wire CLOCK_sgo__sro_n47286;
wire slo__sro_n20322;
wire n_6_2173;
wire n_6_1_280;
wire n_6_2174;
wire n_6_1_281;
wire CLOCK_sgo__n46945;
wire slo__sro_n6229;
wire n_6_2176;
wire slo__sro_n34792;
wire n_6_2177;
wire slo__sro_n29364;
wire n_6_2178;
wire slo__n38401;
wire n_6_2179;
wire n_6_1_286;
wire n_6_2180;
wire slo__sro_n13473;
wire n_6_2181;
wire n_6_1_288;
wire n_6_2182;
wire CLOCK_slo__sro_n50130;
wire n_6_2183;
wire slo__sro_n19568;
wire n_6_2184;
wire slo__n12818;
wire n_6_2185;
wire CLOCK_slo__sro_n50300;
wire n_6_2186;
wire n_6_1_293;
wire n_6_2187;
wire n_6_1_294;
wire CLOCK_sgo__sro_n47262;
wire n_6_1_295;
wire n_6_2189;
wire CLOCK_sgo__sro_n47371;
wire n_6_2190;
wire slo__sro_n13355;
wire n_6_2191;
wire slo__sro_n6160;
wire n_6_2192;
wire slo__sro_n4176;
wire n_6_2193;
wire slo__sro_n31050;
wire CLOCK_sgo__sro_n47210;
wire slo__sro_n15668;
wire n_6_2195;
wire CLOCK_slo__sro_n48813;
wire n_6_2196;
wire slo__sro_n28420;
wire n_6_2197;
wire CLOCK_slo__sro_n51092;
wire n_6_2198;
wire n_6_1_305;
wire n_6_2199;
wire n_6_1_306;
wire n_6_1_307;
wire n_6_1_308;
wire n_6_1_309;
wire n_6_1_310;
wire n_6_2200;
wire n_6_1_311;
wire CLOCK_sgo__sro_n47664;
wire CLOCK_slo__sro_n59641;
wire n_6_2202;
wire slo__n38665;
wire n_6_2203;
wire n_6_1_314;
wire n_6_2204;
wire slo__n41748;
wire n_6_2205;
wire slo__sro_n6654;
wire n_6_2206;
wire slo__n39714;
wire n_6_2207;
wire slo__sro_n12328;
wire n_6_2208;
wire slo__sro_n23159;
wire n_6_2209;
wire n_6_1_320;
wire n_6_2210;
wire slo__sro_n5118;
wire n_6_2211;
wire CLOCK_slo__sro_n50096;
wire n_6_2212;
wire slo__sro_n3905;
wire n_6_2213;
wire n_6_1_324;
wire n_6_2214;
wire n_6_1_325;
wire n_6_2215;
wire slo__sro_n6869;
wire n_6_2216;
wire slo__sro_n36478;
wire n_6_2217;
wire n_6_1_328;
wire slo__sro_n37541;
wire n_6_1_329;
wire n_6_2219;
wire n_6_1_330;
wire n_6_2220;
wire slo__n4932;
wire n_6_2221;
wire slo__sro_n19695;
wire n_6_2222;
wire slo__sro_n9242;
wire n_6_2223;
wire slo__sro_n9815;
wire n_6_2224;
wire n_6_1_335;
wire n_6_2225;
wire slo__n15804;
wire slo__sro_n3056;
wire slo__sro_n19776;
wire n_6_2228;
wire slo__sro_n9845;
wire n_6_2229;
wire n_6_1_340;
wire n_6_2230;
wire n_6_1_341;
wire n_6_1_342;
wire n_6_1_343;
wire n_6_1_344;
wire n_6_1_345;
wire n_6_2231;
wire n_6_1_346;
wire n_6_2232;
wire n_6_1_347;
wire n_6_2233;
wire slo__sro_n9341;
wire n_6_2234;
wire n_6_1_349;
wire n_6_2235;
wire slo__sro_n9343;
wire n_6_2236;
wire slo__sro_n5965;
wire n_6_2237;
wire CLOCK_slo__sro_n49772;
wire n_6_2238;
wire slo__sro_n20260;
wire CLOCK_slo__sro_n48635;
wire n_6_1_354;
wire n_6_2240;
wire slo__sro_n28592;
wire n_6_2241;
wire n_6_1_356;
wire n_6_2242;
wire n_6_1_357;
wire n_6_2243;
wire n_6_1_358;
wire n_6_2244;
wire n_6_1_359;
wire n_6_2245;
wire CLOCK_slo__sro_n48958;
wire n_6_2246;
wire n_6_1_361;
wire n_6_2247;
wire slo__n35483;
wire n_6_2248;
wire slo__sro_n32117;
wire n_6_2249;
wire n_6_1_364;
wire n_6_2250;
wire n_6_1_365;
wire slo__sro_n32317;
wire CLOCK_slo__sro_n53405;
wire n_6_2252;
wire slo__sro_n38699;
wire n_6_2253;
wire n_6_1_368;
wire n_6_2254;
wire n_6_1_369;
wire n_6_2255;
wire slo__sro_n39379;
wire n_6_2256;
wire n_6_1_371;
wire n_6_2257;
wire slo__sro_n9559;
wire n_6_2258;
wire slo__sro_n5056;
wire n_6_2259;
wire slo__sro_n9948;
wire n_6_2260;
wire n_6_1_375;
wire n_6_2261;
wire n_6_1_376;
wire n_6_1_377;
wire n_6_1_378;
wire n_6_1_379;
wire n_6_1_380;
wire n_6_2262;
wire n_6_1_381;
wire n_6_2263;
wire CLOCK_slo__n56284;
wire slo__sro_n6689;
wire CLOCK_sgo__sro_n47732;
wire n_6_1_384;
wire n_6_2266;
wire slo__sro_n9342;
wire n_6_2267;
wire slo__sro_n29674;
wire n_6_2268;
wire slo__sro_n6673;
wire n_6_2269;
wire slo__sro_n6241;
wire n_6_2270;
wire slo__sro_n9671;
wire n_6_2271;
wire slo__n31336;
wire slo__sro_n28562;
wire n_6_2273;
wire slo__sro_n11436;
wire n_6_2274;
wire CLOCK_slo__sro_n59342;
wire n_6_2275;
wire n_6_1_394;
wire slo__sro_n6827;
wire n_6_2277;
wire n_6_1_396;
wire n_6_2278;
wire n_6_1_397;
wire n_6_1_398;
wire n_6_2280;
wire slo__sro_n31087;
wire n_6_2281;
wire slo__sro_n14081;
wire slo__n37549;
wire slo__sro_n19436;
wire n_6_2283;
wire CLOCK_sgo__n48020;
wire n_6_2284;
wire slo__sro_n33595;
wire n_6_2285;
wire slo__sro_n6088;
wire n_6_2286;
wire slo__sro_n12647;
wire n_6_2287;
wire slo__sro_n11796;
wire slo__sro_n19696;
wire n_6_2289;
wire slo__sro_n10458;
wire slo__sro_n28591;
wire slo__sro_n11641;
wire n_6_2291;
wire CLOCK_slo__sro_n54056;
wire n_6_2292;
wire n_6_1_411;
wire n_6_1_412;
wire n_6_1_413;
wire n_6_1_414;
wire n_6_1_415;
wire n_6_2293;
wire slo__sro_n22431;
wire n_6_2294;
wire slo__n18079;
wire n_6_2295;
wire slo__sro_n5875;
wire CLOCK_sgo__sro_n47370;
wire n_6_1_419;
wire n_6_2297;
wire CLOCK_slo__sro_n51723;
wire n_6_2298;
wire n_6_2299;
wire slo__sro_n12225;
wire n_6_2300;
wire slo__n17720;
wire n_6_2301;
wire slo__sro_n9712;
wire n_6_2302;
wire slo__sro_n9701;
wire n_6_2303;
wire slo__sro_n20066;
wire n_6_2304;
wire slo__sro_n40962;
wire n_6_2305;
wire slo__sro_n6897;
wire n_6_2306;
wire slo__sro_n16936;
wire n_6_2307;
wire slo__sro_n21662;
wire n_6_2308;
wire slo__n39180;
wire n_6_2309;
wire slo__sro_n4338;
wire n_6_2310;
wire n_6_1_433;
wire n_6_2311;
wire n_6_1_434;
wire n_6_2312;
wire CLOCK_slo__sro_n52634;
wire n_6_2313;
wire n_6_1_436;
wire n_6_2314;
wire slo__sro_n6367;
wire n_6_2315;
wire n_6_1_438;
wire n_6_2316;
wire n_6_1_439;
wire n_6_2317;
wire n_6_1_440;
wire n_6_2318;
wire slo__sro_n6652;
wire n_6_2319;
wire n_6_1_442;
wire n_6_2320;
wire slo__n12014;
wire slo__sro_n40460;
wire n_6_1_444;
wire n_6_2322;
wire n_6_1_445;
wire n_6_2323;
wire n_6_1_446;
wire n_6_1_447;
wire n_6_1_448;
wire n_6_1_449;
wire n_6_1_450;
wire n_6_2324;
wire n_6_1_451;
wire CLOCK_sgo__sro_n47760;
wire n_6_1_452;
wire slo__sro_n30705;
wire slo__sro_n6829;
wire slo__sro_n30363;
wire n_6_1_454;
wire drc_ipo_n26606;
wire slo__n29454;
wire n_6_2329;
wire n_6_1_456;
wire n_6_2330;
wire n_6_1_457;
wire drc_ipo_n26599;
wire n_6_1_458;
wire slo__sro_n36477;
wire n_6_2333;
wire slo__n11420;
wire n_6_2334;
wire slo__sro_n7186;
wire n_6_2335;
wire slo__sro_n16920;
wire n_6_2336;
wire slo___n17155;
wire n_6_2337;
wire n_6_1_464;
wire n_6_2338;
wire slo__sro_n5711;
wire n_6_2339;
wire slo__sro_n8918;
wire n_6_2340;
wire CLOCK_slo__sro_n52670;
wire n_6_2341;
wire slo__sro_n10270;
wire n_6_2342;
wire n_6_1_469;
wire n_6_2343;
wire n_6_1_470;
wire n_6_2344;
wire n_6_2345;
wire slo__n17435;
wire n_6_2346;
wire slo__sro_n19805;
wire slo__sro_n32319;
wire slo__sro_n28419;
wire n_6_2348;
wire n_6_1_475;
wire n_6_2349;
wire slo__sro_n17753;
wire n_6_2350;
wire slo__sro_n38744;
wire n_6_2351;
wire spt__n66402;
wire n_6_2352;
wire n_6_1_479;
wire CLOCK_sgo__sro_n47287;
wire CLOCK_slo__sro_n52136;
wire n_6_2354;
wire n_6_1_481;
wire n_6_1_482;
wire n_6_1_483;
wire n_6_1_484;
wire n_6_1_485;
wire n_6_2355;
wire n_6_1_486;
wire n_6_2356;
wire n_6_1_487;
wire n_6_2357;
wire n_6_1_488;
wire slo__sro_n31051;
wire n_6_1_489;
wire n_6_2359;
wire slo__n17338;
wire n_6_2360;
wire slo__sro_n32138;
wire n_6_2361;
wire n_6_1_492;
wire n_6_2362;
wire slo__sro_n20885;
wire drc_ipo_n26601;
wire n_6_2364;
wire CLOCK_slo__sro_n52916;
wire n_6_2365;
wire n_6_1_496;
wire n_6_2366;
wire slo__n30671;
wire n_6_2367;
wire slo__sro_n20394;
wire n_6_2368;
wire slo__sro_n5877;
wire drc_ipo_n26605;
wire slo__sro_n34276;
wire n_6_2370;
wire n_6_1_501;
wire n_6_2371;
wire slo__sro_n5855;
wire n_6_2372;
wire CLOCK_slo__sro_n61308;
wire n_6_2373;
wire n_6_1_504;
wire n_6_2374;
wire n_6_1_505;
wire n_6_2375;
wire CLOCK_slo__sro_n51979;
wire n_6_2376;
wire n_6_1_507;
wire n_6_2377;
wire slo__sro_n4784;
wire n_6_2378;
wire n_6_1_509;
wire n_6_2379;
wire slo__sro_n27836;
wire n_6_2380;
wire n_6_1_511;
wire n_6_2381;
wire slo__n17713;
wire n_6_2382;
wire n_6_1_513;
wire n_6_2383;
wire n_6_1_514;
wire n_6_2384;
wire n_6_1_515;
wire CLOCK_sgo__sro_n47297;
wire n_6_1_516;
wire n_6_1_517;
wire n_6_1_518;
wire n_6_1_519;
wire n_6_1_520;
wire n_6_2386;
wire n_6_1_521;
wire slo__sro_n30995;
wire n_6_1_522;
wire n_6_2388;
wire n_6_1_523;
wire CLOCK_slo__n64837;
wire n_6_1_524;
wire n_6_2390;
wire slo__sro_n6870;
wire n_6_2391;
wire n_6_1_526;
wire n_6_2392;
wire slo__sro_n7690;
wire n_6_2393;
wire n_6_1_528;
wire n_6_2394;
wire slo__n36610;
wire n_6_2395;
wire slo__sro_n7371;
wire CLOCK_slo__sro_n55059;
wire slo__sro_n41479;
wire n_6_2397;
wire n_6_1_532;
wire n_6_2398;
wire slo__sro_n7833;
wire slo__sro_n35184;
wire slo__sro_n33562;
wire n_6_2401;
wire n_6_1_536;
wire n_6_2402;
wire CLOCK_slo__sro_n54101;
wire n_6_2403;
wire CLOCK_slo__n64621;
wire n_6_2404;
wire n_6_1_539;
wire n_6_2405;
wire n_6_1_540;
wire n_6_2406;
wire slo__sro_n31817;
wire slo__sro_n42343;
wire n_6_1_542;
wire n_6_2408;
wire slo__sro_n8171;
wire n_6_2409;
wire slo__sro_n4814;
wire n_6_2410;
wire n_6_1_545;
wire n_6_2411;
wire slo__sro_n19806;
wire n_6_2412;
wire n_6_1_547;
wire n_6_2413;
wire n_6_1_548;
wire n_6_2414;
wire n_6_1_549;
wire n_6_2415;
wire n_6_1_550;
wire n_6_2416;
wire slo__sro_n36849;
wire n_6_1_552;
wire n_6_1_553;
wire n_6_1_554;
wire n_6_1_555;
wire n_6_2417;
wire n_6_1_556;
wire n_6_2418;
wire n_6_1_557;
wire n_6_2419;
wire slo__sro_n7306;
wire n_6_2420;
wire slo__sro_n7270;
wire n_6_2421;
wire slo__sro_n7435;
wire n_6_2422;
wire slo__sro_n7772;
wire n_6_2423;
wire n_6_1_562;
wire n_6_2424;
wire n_6_1_563;
wire n_6_2425;
wire slo__n28538;
wire n_6_2426;
wire slo__sro_n28006;
wire CLOCK_slo__sro_n51595;
wire CLOCK_slo__sro_n65030;
wire CLOCK_slo__sro_n48815;
wire n_6_1_567;
wire n_6_2429;
wire slo__sro_n19997;
wire n_6_2430;
wire slo__sro_n19973;
wire n_6_2431;
wire slo__mro_n33047;
wire n_6_2432;
wire n_6_1_571;
wire n_6_2433;
wire n_6_1_572;
wire slo__sro_n10427;
wire n_6_2435;
wire n_6_1_574;
wire n_6_2436;
wire n_6_1_575;
wire n_6_2437;
wire CLOCK_slo__sro_n59467;
wire n_6_2438;
wire n_6_1_577;
wire n_6_2439;
wire slo__sro_n33597;
wire n_6_2440;
wire slo__sro_n33777;
wire slo__sro_n37974;
wire n_6_1_580;
wire n_6_2442;
wire n_6_1_581;
wire slo__sro_n29443;
wire slo__sro_n21795;
wire n_6_2444;
wire slo__sro_n33788;
wire slo__sro_n40770;
wire CLOCK_slo__sro_n55102;
wire n_6_2446;
wire n_6_1_585;
wire n_6_2447;
wire n_6_1_586;
wire n_6_1_587;
wire n_6_1_588;
wire n_6_1_589;
wire n_6_1_590;
wire n_6_2448;
wire n_6_1_591;
wire slo__sro_n31656;
wire n_6_1_592;
wire n_6_2450;
wire n_6_1_593;
wire n_6_2451;
wire slo__sro_n7466;
wire n_6_2452;
wire n_6_1_595;
wire n_6_2453;
wire slo__sro_n21676;
wire drc_ipo_n26600;
wire slo__sro_n20613;
wire n_6_2455;
wire slo__sro_n20734;
wire n_6_2456;
wire CLOCK_slo__sro_n50658;
wire n_6_2457;
wire n_6_1_600;
wire opt_ipo_n45565;
wire n_6_1_601;
wire n_6_2459;
wire n_6_1_602;
wire n_6_2460;
wire slo__sro_n36476;
wire n_6_2461;
wire n_6_1_604;
wire n_6_2462;
wire slo__sro_n28681;
wire n_6_2463;
wire slo__sro_n37819;
wire n_6_2464;
wire slo__sro_n20321;
wire n_6_2465;
wire slo__n14148;
wire n_6_2466;
wire CLOCK_slo__sro_n59437;
wire n_6_2467;
wire CLOCK_slo__sro_n51511;
wire n_6_2468;
wire n_6_1_611;
wire n_6_2469;
wire slo__sro_n19752;
wire n_6_2470;
wire n_6_1_613;
wire n_6_2471;
wire CLOCK_slo__sro_n51541;
wire n_6_2472;
wire slo__sro_n5865;
wire n_6_1_616;
wire n_6_2474;
wire slo__sro_n12506;
wire n_6_2475;
wire n_6_2476;
wire slo__sro_n20923;
wire n_6_2477;
wire n_6_1_620;
wire n_6_2478;
wire n_6_1_621;
wire n_6_1_622;
wire n_6_1_623;
wire n_6_1_624;
wire n_6_1_625;
wire n_6_2479;
wire n_6_1_626;
wire n_6_2480;
wire n_6_1_627;
wire n_6_2481;
wire slo__sro_n21632;
wire n_6_2482;
wire n_6_1_629;
wire n_6_2483;
wire n_6_1_630;
wire n_6_2484;
wire slo__sro_n9122;
wire n_6_2485;
wire n_6_1_632;
wire n_6_2486;
wire slo__n17556;
wire n_6_2487;
wire n_6_1_634;
wire n_6_2488;
wire n_6_1_635;
wire n_6_2489;
wire CLOCK_slo__sro_n51261;
wire n_6_2490;
wire slo__sro_n34279;
wire n_6_2491;
wire slo__sro_n4529;
wire n_6_2492;
wire n_6_1_639;
wire n_6_2493;
wire CLOCK_slo__sro_n62841;
wire n_6_2494;
wire slo__n14603;
wire n_6_2495;
wire slo__sro_n38758;
wire n_6_2496;
wire slo__sro_n21437;
wire n_6_2497;
wire n_6_1_644;
wire n_6_2498;
wire n_6_1_645;
wire n_6_2499;
wire n_6_1_646;
wire n_6_2500;
wire slo__mro_n33032;
wire n_6_2501;
wire n_6_1_648;
wire n_6_2502;
wire n_6_1_649;
wire n_6_2503;
wire n_6_1_650;
wire n_6_2504;
wire slo__sro_n7692;
wire n_6_2505;
wire n_6_1_652;
wire n_6_2506;
wire CLOCK_slo__sro_n50318;
wire n_6_2507;
wire spw__n67541;
wire n_6_2508;
wire n_6_1_655;
wire n_6_2509;
wire n_6_1_656;
wire n_6_1_657;
wire n_6_1_658;
wire n_6_1_659;
wire n_6_1_660;
wire n_6_2510;
wire n_6_1_661;
wire n_6_2511;
wire CLOCK_slo__sro_n49402;
wire slo__sro_n30997;
wire slo__sro_n7583;
wire n_6_2513;
wire CLOCK_slo__sro_n60762;
wire n_6_2514;
wire slo__sro_n31219;
wire drc_ipo_n26596;
wire slo__sro_n9138;
wire drc_ipo_n26597;
wire n_6_1_667;
wire n_6_2517;
wire slo__sro_n36945;
wire n_6_2518;
wire n_6_1_669;
wire n_6_2519;
wire n_6_1_670;
wire n_6_2520;
wire slo__sro_n34554;
wire CLOCK_slo__sro_n61283;
wire slo__n32747;
wire opt_ipo_n23778;
wire slo__sro_n7705;
wire n_6_2523;
wire slo__sro_n7405;
wire n_6_2524;
wire n_6_1_675;
wire n_6_2525;
wire n_6_1_676;
wire n_6_2526;
wire slo__sro_n30032;
wire n_6_2527;
wire slo__sro_n7910;
wire n_6_2528;
wire slo__sro_n9268;
wire n_6_2529;
wire CLOCK_slo__sro_n54647;
wire n_6_2530;
wire CLOCK_slo__sro_n53420;
wire n_6_2531;
wire n_6_1_682;
wire n_6_2532;
wire slo__sro_n8684;
wire n_6_2533;
wire n_6_1_684;
wire n_6_2534;
wire n_6_1_685;
wire n_6_2535;
wire slo__sro_n30146;
wire drc_ipo_n26602;
wire n_6_1_687;
wire n_6_2537;
wire CLOCK_slo__n55287;
wire n_6_2538;
wire CLOCK_slo__sro_n55168;
wire n_6_2539;
wire n_6_1_690;
wire n_6_2540;
wire n_6_1_691;
wire n_6_1_692;
wire n_6_1_693;
wire n_6_1_694;
wire n_6_1_695;
wire n_6_2541;
wire n_6_1_696;
wire n_6_2542;
wire n_6_1_697;
wire n_6_2543;
wire CLOCK_slo__sro_n63005;
wire n_6_2544;
wire n_6_1_699;
wire n_6_2545;
wire n_6_1_700;
wire n_6_2546;
wire slo__sro_n12410;
wire n_6_2547;
wire slo__sro_n42341;
wire n_6_2548;
wire n_6_1_703;
wire n_6_2549;
wire n_6_1_704;
wire spw__n68268;
wire slo__sro_n14857;
wire n_6_2551;
wire n_6_1_706;
wire n_6_2552;
wire n_6_1_707;
wire n_6_2553;
wire n_6_2554;
wire slo__n14899;
wire n_6_2555;
wire slo__sro_n8179;
wire n_6_2556;
wire n_6_1_711;
wire n_6_2557;
wire n_6_1_712;
wire n_6_2558;
wire n_6_1_713;
wire n_6_2559;
wire n_6_1_714;
wire n_6_2560;
wire slo__sro_n12490;
wire n_6_2561;
wire slo__sro_n33790;
wire n_6_2562;
wire n_6_1_717;
wire n_6_2563;
wire n_6_1_718;
wire n_6_2564;
wire n_6_1_719;
wire n_6_2565;
wire n_6_1_720;
wire n_6_2566;
wire slo__sro_n32203;
wire n_6_2567;
wire slo__sro_n10098;
wire n_6_2568;
wire n_6_1_723;
wire n_6_2569;
wire n_6_1_724;
wire n_6_2570;
wire n_6_1_725;
wire n_6_2571;
wire n_6_1_726;
wire n_6_1_727;
wire n_6_1_728;
wire n_6_1_729;
wire n_6_1_730;
wire n_6_2572;
wire n_6_1_731;
wire n_6_2573;
wire n_6_1_732;
wire n_6_2574;
wire n_6_1_733;
wire CLOCK_slo__sro_n49243;
wire n_6_1_734;
wire n_6_2576;
wire slo__sro_n11474;
wire n_6_2577;
wire slo__sro_n35183;
wire CLOCK_opt_ipo_n46124;
wire slo__sro_n14854;
wire drc_ipo_n26592;
wire slo___n7881;
wire CLOCK_slo__sro_n48977;
wire slo__sro_n37192;
wire n_6_2581;
wire slo__sro_n27689;
wire n_6_2582;
wire n_6_1_741;
wire n_6_2583;
wire slo__n14942;
wire n_6_2584;
wire n_6_1_743;
wire n_6_2585;
wire n_6_1_744;
wire n_6_2586;
wire n_6_1_745;
wire n_6_2587;
wire slo__sro_n10271;
wire n_6_2588;
wire CLOCK_slo__sro_n51132;
wire n_6_2589;
wire n_6_1_748;
wire n_6_2590;
wire n_6_1_749;
wire n_6_2591;
wire CLOCK_slo__sro_n55929;
wire n_6_2592;
wire slo__sro_n29017;
wire n_6_2593;
wire slo__sro_n35197;
wire n_6_2594;
wire slo__sro_n22132;
wire n_6_2595;
wire n_6_1_754;
wire n_6_2596;
wire n_6_1_755;
wire n_6_2597;
wire n_6_1_756;
wire slo__sro_n29653;
wire n_6_1_757;
wire slo__n35802;
wire CLOCK_slo__sro_n65090;
wire n_6_2600;
wire n_6_1_759;
wire n_6_2601;
wire n_6_1_760;
wire n_6_2602;
wire n_6_1_761;
wire n_6_1_762;
wire n_6_1_763;
wire n_6_1_764;
wire n_6_1_765;
wire spc__n66318;
wire n_6_1_766;
wire n_6_2604;
wire n_6_1_767;
wire CLOCK_slo__sro_n62895;
wire slo__sro_n41061;
wire CLOCK_slo__sro_n58343;
wire n_6_2607;
wire n_6_1_770;
wire n_6_2608;
wire slo__sro_n34553;
wire n_6_2609;
wire slo__sro_n5678;
wire n_6_2610;
wire n_6_1_773;
wire n_6_2611;
wire slo__sro_n32044;
wire n_6_2612;
wire n_6_1_775;
wire n_6_2613;
wire slo__sro_n10378;
wire n_6_2614;
wire n_6_1_777;
wire n_6_2615;
wire slo__sro_n16216;
wire n_6_2616;
wire n_6_1_779;
wire n_6_2617;
wire CLOCK_slo__sro_n49242;
wire n_6_2618;
wire CLOCK_slo__sro_n51765;
wire drc_ipo_n26595;
wire n_6_1_782;
wire slo__sro_n29774;
wire slo___n13099;
wire n_6_2621;
wire slo__sro_n6651;
wire n_6_2622;
wire slo__n19260;
wire n_6_2623;
wire slo__sro_n7944;
wire drc_ipo_n26598;
wire slo__n12976;
wire n_6_2625;
wire n_6_1_788;
wire n_6_2626;
wire n_6_1_789;
wire n_6_2627;
wire n_6_1_790;
wire n_6_2628;
wire n_6_1_791;
wire n_6_2629;
wire n_6_1_792;
wire n_6_2630;
wire n_6_1_793;
wire n_6_2631;
wire n_6_1_794;
wire n_6_2632;
wire n_6_1_795;
wire n_6_2633;
wire n_6_1_796;
wire n_6_1_797;
wire n_6_1_798;
wire n_6_1_799;
wire n_6_1_800;
wire n_6_2634;
wire n_6_1_801;
wire n_6_2635;
wire n_6_1_802;
wire n_6_2636;
wire n_6_1_803;
wire n_6_2637;
wire slo__sro_n35185;
wire n_6_2638;
wire CLOCK_slo__sro_n48698;
wire n_6_2639;
wire n_6_1_806;
wire n_6_2640;
wire slo__sro_n29880;
wire n_6_2641;
wire n_6_1_808;
wire n_6_2642;
wire n_6_1_809;
wire drc_ipo_n26591;
wire slo__sro_n6239;
wire n_6_2644;
wire n_6_1_811;
wire n_6_2645;
wire CLOCK_slo__sro_n53080;
wire n_6_2646;
wire n_6_1_813;
wire n_6_2647;
wire slo__sro_n7423;
wire n_6_2648;
wire n_6_1_815;
wire n_6_2649;
wire CLOCK_slo__sro_n63268;
wire n_6_2650;
wire n_6_2651;
wire slo__sro_n19970;
wire n_6_2652;
wire n_6_1_819;
wire n_6_2653;
wire n_6_1_820;
wire CLOCK_slo__sro_n62823;
wire slo__sro_n8580;
wire drc_ipo_n26594;
wire slo__sro_n8602;
wire n_6_2656;
wire CLOCK_slo__sro_n56596;
wire n_6_2657;
wire n_6_1_824;
wire n_6_2658;
wire n_6_1_825;
wire n_6_2659;
wire slo__n11409;
wire n_6_2660;
wire n_6_1_827;
wire n_6_2661;
wire n_6_1_828;
wire n_6_2662;
wire n_6_1_829;
wire n_6_2663;
wire n_6_1_830;
wire n_6_2664;
wire n_6_1_831;
wire n_6_1_832;
wire CLOCK_slo__sro_n61347;
wire n_6_1_834;
wire n_6_1_835;
wire n_6_2665;
wire n_6_1_836;
wire n_6_2666;
wire slo__sro_n7406;
wire n_6_2667;
wire slo__sro_n4774;
wire n_6_2668;
wire n_6_1_839;
wire CLOCK_slo__n48588;
wire slo__sro_n15199;
wire n_6_2670;
wire slo___n19058;
wire CLOCK_slo__sro_n48634;
wire slo__sro_n6791;
wire n_6_2672;
wire slo__sro_n7912;
wire n_6_2673;
wire CLOCK_sgo__sro_n47369;
wire CLOCK_slo__sro_n62332;
wire slo__sro_n8777;
wire n_6_2675;
wire slo__sro_n34136;
wire n_6_2676;
wire slo__sro_n34277;
wire n_6_2677;
wire slo__n35733;
wire n_6_2678;
wire n_6_1_849;
wire n_6_2679;
wire slo__sro_n37539;
wire n_6_2680;
wire n_6_1_851;
wire n_6_2681;
wire CLOCK_slo__sro_n49603;
wire n_6_2682;
wire slo__sro_n37209;
wire n_6_2683;
wire slo__sro_n8582;
wire n_6_2684;
wire slo__sro_n19960;
wire n_6_2685;
wire slo__sro_n7617;
wire n_6_2686;
wire n_6_1_857;
wire slo__sro_n26912;
wire spw__n67889;
wire n_6_2688;
wire slo__sro_n8310;
wire n_6_2689;
wire slo___n9717;
wire n_6_2690;
wire n_6_1_861;
wire CLOCK_sgo__sro_n47801;
wire n_6_1_862;
wire n_6_2692;
wire slo__sro_n4286;
wire n_6_2693;
wire n_6_1_864;
wire n_6_2694;
wire n_6_1_865;
wire n_6_2695;
wire n_6_1_866;
wire n_6_1_867;
wire n_6_1_868;
wire n_6_1_869;
wire n_6_1_870;
wire n_6_2696;
wire n_6_1_871;
wire slo__mro_n32529;
wire CLOCK_slo__sro_n63090;
wire n_6_2698;
wire n_6_1_873;
wire CLOCK_sgo__sro_n47244;
wire n_6_1_874;
wire CLOCK_slo__sro_n49385;
wire n_6_1_875;
wire n_6_2701;
wire slo__sro_n31830;
wire n_6_2702;
wire n_6_1_877;
wire n_6_2703;
wire n_6_1_878;
wire n_6_2704;
wire n_6_1_879;
wire slo__sro_n29859;
wire n_6_1_880;
wire drc_ipo_n26589;
wire n_6_1_881;
wire n_6_2707;
wire n_6_1_882;
wire drc_ipo_n26590;
wire n_6_1_883;
wire n_6_2709;
wire n_6_1_884;
wire n_6_2710;
wire n_6_1_885;
wire n_6_2711;
wire n_6_1_886;
wire n_6_2712;
wire n_6_1_887;
wire n_6_2713;
wire n_6_1_888;
wire n_6_2714;
wire slo__n13938;
wire n_6_2715;
wire slo__sro_n37389;
wire n_6_2716;
wire n_6_1_891;
wire n_6_2717;
wire n_6_1_892;
wire n_6_2718;
wire CLOCK_slo__sro_n56894;
wire n_6_2719;
wire n_6_1_894;
wire n_6_2720;
wire slo__sro_n8834;
wire n_6_2721;
wire slo__sro_n8978;
wire n_6_2722;
wire slo__sro_n34620;
wire n_6_2723;
wire n_6_1_898;
wire n_6_2724;
wire slo__n30795;
wire n_6_2725;
wire n_6_1_900;
wire n_6_2726;
wire n_6_1_901;
wire n_6_1_902;
wire CLOCK_slo__sro_n61295;
wire n_6_1_904;
wire n_6_1_905;
wire n_6_2727;
wire n_6_1_906;
wire n_6_2728;
wire n_6_1_907;
wire n_6_2729;
wire slo___n8281;
wire n_6_2730;
wire n_6_1_909;
wire n_6_2731;
wire slo__sro_n7945;
wire n_6_2732;
wire n_6_1_911;
wire CLOCK_sgo__sro_n47561;
wire slo__n14696;
wire CLOCK_opt_ipo_n45893;
wire slo__sro_n8339;
wire n_6_2735;
wire slo__sro_n15185;
wire n_6_2736;
wire n_6_1_915;
wire n_6_2737;
wire slo__sro_n9421;
wire n_6_2738;
wire n_6_1_917;
wire n_6_2739;
wire slo__sro_n12409;
wire n_6_2740;
wire n_6_1_919;
wire n_6_2741;
wire n_6_1_920;
wire n_6_2742;
wire slo__sro_n5416;
wire n_6_2743;
wire slo__sro_n22702;
wire n_6_2744;
wire n_6_1_923;
wire n_6_2745;
wire slo__sro_n9561;
wire n_6_2746;
wire n_6_1_925;
wire n_6_2747;
wire n_6_1_926;
wire n_6_2748;
wire n_6_1_927;
wire n_6_2749;
wire slo__sro_n11858;
wire n_6_2750;
wire n_6_1_929;
wire n_6_2751;
wire n_6_1_930;
wire n_6_2752;
wire n_6_1_931;
wire opt_ipo_n45324;
wire slo__sro_n8991;
wire n_6_2754;
wire n_6_1_933;
wire n_6_2755;
wire CLOCK_slo__sro_n59729;
wire n_6_2756;
wire n_6_1_935;
wire n_6_2757;
wire n_6_1_936;
wire n_6_1_937;
wire CLOCK_slo__sro_n61783;
wire n_6_1_939;
wire n_6_1_940;
wire n_6_2758;
wire n_6_1_941;
wire n_6_2759;
wire n_6_1_942;
wire n_6_2760;
wire n_6_1_943;
wire slo__sro_n31361;
wire slo__sro_n27860;
wire n_6_2762;
wire n_6_1_945;
wire n_6_2763;
wire n_6_1_946;
wire CLOCK_slo__n48618;
wire slo__sro_n35186;
wire CLOCK_slo__sro_n56608;
wire slo__sro_n8900;
wire n_6_2766;
wire n_6_1_949;
wire n_6_2767;
wire n_6_1_950;
wire n_6_2768;
wire n_6_1_951;
wire n_6_2769;
wire slo__n10924;
wire n_6_2770;
wire slo__n11048;
wire n_6_2771;
wire CLOCK_opt_ipo_n45744;
wire n_6_2772;
wire slo__sro_n10272;
wire n_6_2773;
wire n_6_1_956;
wire n_6_2774;
wire slo__sro_n9533;
wire n_6_2775;
wire CLOCK_slo__sro_n59304;
wire n_6_2776;
wire slo__sro_n27581;
wire n_6_2777;
wire n_6_1_960;
wire n_6_2778;
wire slo__sro_n36683;
wire n_6_2779;
wire n_6_1_962;
wire n_6_2780;
wire CLOCK_sgo__sro_n48085;
wire n_6_2781;
wire slo__sro_n15108;
wire n_6_2782;
wire n_6_1_965;
wire CLOCK_slo__sro_n49673;
wire n_6_1_966;
wire n_6_2784;
wire n_6_1_967;
wire n_6_2785;
wire n_6_1_968;
wire n_6_2786;
wire n_6_1_969;
wire n_6_2787;
wire n_6_1_970;
wire n_6_2788;
wire n_6_1_971;
wire n_6_1_972;
wire n_6_1_973;
wire n_6_1_974;
wire n_6_1_975;
wire n_6_2789;
wire n_6_1_976;
wire n_6_2790;
wire CLOCK_slo__sro_n64180;
wire n_6_2791;
wire slo__sro_n20666;
wire n_6_2792;
wire n_6_1_979;
wire n_6_2793;
wire slo___n23215;
wire n_6_2794;
wire slo__sro_n33776;
wire n_6_2795;
wire slo__sro_n35270;
wire n_6_2796;
wire n_6_1_983;
wire CLOCK_slo__sro_n62668;
wire n_6_1_984;
wire CLOCK_sgo__sro_n47665;
wire n_6_1_985;
wire n_6_2799;
wire slo__sro_n32027;
wire n_6_2800;
wire slo__sro_n35509;
wire n_6_2801;
wire slo__n18286;
wire n_6_2802;
wire CLOCK_slo__sro_n62489;
wire n_6_2803;
wire CLOCK_slo__sro_n65088;
wire n_6_2804;
wire n_6_1_991;
wire n_6_2805;
wire n_6_1_992;
wire slo__sro_n34757;
wire n_6_1_993;
wire n_6_2807;
wire n_6_1_994;
wire CLOCK_slo__sro_n50792;
wire n_6_1_995;
wire n_6_2809;
wire CLOCK_slo__n56075;
wire n_6_2810;
wire slo__n14062;
wire n_6_2811;
wire n_6_1_998;
wire n_6_2812;
wire slo__sro_n11594;
wire n_6_2813;
wire n_6_1_1000;
wire drc_ipo_n26588;
wire n_6_1_1001;
wire n_6_2815;
wire slo__sro_n11844;
wire n_6_2816;
wire slo__sro_n12110;
wire n_6_2817;
wire n_6_1_1004;
wire n_6_2818;
wire slo__sro_n22735;
wire n_6_1_1006;
wire n_6_1_1007;
wire CLOCK_slo__sro_n61349;
wire n_6_1_1009;
wire n_6_1_1010;
wire n_6_2820;
wire slo__sro_n33706;
wire n_6_2821;
wire CLOCK_slo__sro_n61696;
wire drc_ipo_n26582;
wire slo__sro_n8966;
wire slo__sro_n30019;
wire slo__sro_n9430;
wire CLOCK_slo__sro_n49427;
wire slo__sro_n35288;
wire CLOCK_slo__sro_n49602;
wire CLOCK_slo__sro_n55809;
wire n_6_2826;
wire n_6_1_1017;
wire n_6_2827;
wire n_6_1_1018;
wire n_6_2828;
wire CLOCK_sgo__sro_n47149;
wire n_6_2829;
wire n_6_1_1020;
wire n_6_2830;
wire n_6_1_1021;
wire n_6_2831;
wire slo__sro_n11754;
wire n_6_2832;
wire n_6_1_1023;
wire n_6_2833;
wire n_6_1_1024;
wire n_6_2834;
wire slo__sro_n29857;
wire n_6_2835;
wire slo__sro_n32471;
wire n_6_2836;
wire slo__n37202;
wire CLOCK_slo__sro_n62932;
wire slo__sro_n30031;
wire drc_ipo_n26583;
wire n_6_1_1029;
wire n_6_2839;
wire n_6_1_1030;
wire n_6_2840;
wire slo__sro_n29652;
wire drc_ipo_n26585;
wire n_6_1_1032;
wire n_6_2842;
wire CLOCK_slo__sro_n57315;
wire n_6_2843;
wire n_6_1_1034;
wire n_6_2844;
wire n_6_1_1035;
wire n_6_2845;
wire slo__sro_n8390;
wire n_6_2846;
wire n_6_1_1037;
wire n_6_2847;
wire n_6_1_1038;
wire n_6_2848;
wire slo__sro_n40959;
wire n_6_2849;
wire n_6_1_1040;
wire n_6_2850;
wire n_6_1_1041;
wire n_6_1_1042;
wire CLOCK_slo__sro_n61784;
wire n_6_1_1044;
wire n_6_1_1045;
wire n_6_2851;
wire CLOCK_slo__sro_n61307;
wire n_6_2852;
wire n_6_1_1047;
wire n_6_2853;
wire CLOCK_sgo__sro_n47246;
wire n_6_2854;
wire slo__sro_n9085;
wire n_6_2855;
wire spw__n66887;
wire n_6_2856;
wire slo__sro_n9007;
wire n_6_2857;
wire n_6_1_1052;
wire n_6_2858;
wire n_6_1_1053;
wire n_6_2859;
wire n_6_1_1054;
wire n_6_2860;
wire n_6_1_1055;
wire n_6_2861;
wire slo__n36350;
wire n_6_2862;
wire slo__n35792;
wire n_6_2863;
wire slo__sro_n32212;
wire n_6_2864;
wire n_6_1_1059;
wire n_6_2865;
wire slo__sro_n22347;
wire n_6_2866;
wire slo___n17357;
wire n_6_2867;
wire CLOCK_slo__n62554;
wire n_6_2868;
wire slo__sro_n8500;
wire n_6_2869;
wire slo__sro_n8430;
wire n_6_2870;
wire slo__sro_n39899;
wire n_6_2871;
wire n_6_1_1066;
wire n_6_2872;
wire n_6_1_1067;
wire n_6_2873;
wire slo__sro_n20845;
wire slo__n38656;
wire n_6_1_1069;
wire n_6_2875;
wire slo__sro_n7960;
wire n_6_2876;
wire n_6_1_1071;
wire n_6_2877;
wire n_6_1_1072;
wire drc_ipo_n26584;
wire slo__sro_n7852;
wire slo__sro_n13965;
wire n_6_1_1074;
wire n_6_2880;
wire n_6_1_1075;
wire n_6_2881;
wire n_6_1_1076;
wire n_6_1_1077;
wire drc_ipo_n26579;
wire n_6_1_1079;
wire n_6_1_1080;
wire CLOCK_sgo__n47026;
wire n_6_1_1081;
wire n_6_2883;
wire sgo__sro_n1677;
wire n_6_2884;
wire sgo__sro_n1643;
wire n_6_2885;
wire sgo__sro_n1718;
wire n_6_2886;
wire n_6_1_1085;
wire n_6_2887;
wire sgo__sro_n1719;
wire CLOCK_slo__sro_n49605;
wire slo__sro_n2122;
wire n_6_2889;
wire n_6_1_1088;
wire n_6_2890;
wire n_6_1_1089;
wire n_6_2891;
wire n_6_1_1090;
wire n_6_2892;
wire slo__sro_n2206;
wire n_6_2893;
wire slo__sro_n2194;
wire n_6_2894;
wire slo__sro_n2306;
wire n_6_2895;
wire slo__sro_n2220;
wire n_6_2896;
wire n_6_1_1095;
wire n_6_2897;
wire slo__sro_n2272;
wire n_6_2898;
wire n_6_1_1097;
wire n_6_2899;
wire slo__sro_n2242;
wire n_6_2900;
wire slo__sro_n2284;
wire n_6_2901;
wire n_6_1_1100;
wire n_6_2902;
wire slo__sro_n2362;
wire n_6_2903;
wire n_6_1_1102;
wire n_6_2904;
wire n_6_1_1103;
wire n_6_2905;
wire n_6_1_1104;
wire n_6_2906;
wire n_6_1_1105;
wire n_6_2907;
wire n_6_1_1106;
wire n_6_2908;
wire slo__sro_n2400;
wire n_6_2909;
wire drc_ipo_n26581;
wire n_6_2910;
wire n_6_1_1109;
wire slo__sro_n31798;
wire n_6_2911;
wire n_6_1_1111;
wire drc_ipo_n26576;
wire n_6_2912;
wire n_6_1_1113;
wire n_6_1_1114;
wire n_6_2913;
wire n_6_1_1115;
wire n_6_1_1116;
wire n_6_1_1117;
wire n_6_1_1118;
wire n_6_1_1119;
wire n_6_1_1120;
wire n_6_1_1121;
wire n_6_1_1122;
wire n_6_1_1123;
wire n_6_1_1124;
wire n_6_1_1125;
wire n_6_1_1126;
wire n_6_1_1127;
wire n_6_1_1128;
wire n_6_1_1129;
wire n_6_1_1130;
wire n_6_1_1131;
wire n_6_1_1132;
wire n_6_1_1133;
wire n_6_1_1134;
wire n_6_1_1135;
wire n_6_1_1136;
wire n_6_1_1137;
wire n_6_1_1138;
wire n_6_1_1139;
wire n_6_1_1140;
wire n_6_1_1141;
wire n_6_1_1142;
wire n_6_1_1143;
wire n_6_1_1144;
wire n_6_1_1145;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;
wire n_0_10;
wire n_0_11;
wire n_0_12;
wire n_0_13;
wire n_0_14;
wire n_0_15;
wire n_0_16;
wire n_0_17;
wire n_0_18;
wire n_0_19;
wire n_0_20;
wire n_0_21;
wire n_0_22;
wire n_0_23;
wire n_0_24;
wire n_0_25;
wire n_0_26;
wire n_0_27;
wire n_0_28;
wire n_0_29;
wire n_0_30;
wire n_0_31;
wire n_0_32;
wire n_0_33;
wire n_0_34;
wire n_0_35;
wire n_0_36;
wire n_0_37;
wire n_0_38;
wire n_0_39;
wire n_0_40;
wire n_0_41;
wire n_0_42;
wire n_0_43;
wire n_0_44;
wire n_0_45;
wire n_0_46;
wire n_0_47;
wire n_0_48;
wire n_0_49;
wire n_0_50;
wire n_0_51;
wire n_0_52;
wire n_0_53;
wire n_0_54;
wire n_0_55;
wire n_0_56;
wire n_0_57;
wire n_0_58;
wire n_0_59;
wire n_0_60;
wire n_0_61;
wire n_0_62;
wire n_0_0_0;
wire n_0_0_1;
wire n_0_63;
wire n_0_64;
wire n_0_65;
wire n_0_66;
wire n_0_67;
wire n_0_68;
wire n_0_69;
wire n_0_70;
wire n_0_71;
wire n_0_72;
wire n_0_73;
wire n_0_74;
wire n_0_75;
wire n_0_76;
wire n_0_77;
wire n_0_78;
wire n_0_79;
wire n_0_80;
wire n_0_81;
wire n_0_82;
wire n_0_83;
wire n_0_84;
wire n_0_85;
wire n_0_86;
wire n_0_87;
wire n_0_88;
wire n_0_89;
wire n_0_90;
wire n_0_91;
wire n_0_92;
wire n_0_93;
wire n_0_94;
wire n_0_95;
wire n_0_96;
wire n_0_97;
wire n_0_98;
wire n_0_99;
wire n_0_100;
wire n_0_101;
wire n_0_102;
wire n_0_103;
wire n_0_104;
wire n_0_105;
wire n_0_106;
wire n_0_107;
wire n_0_108;
wire n_0_109;
wire n_0_110;
wire n_0_111;
wire n_0_112;
wire n_0_113;
wire n_0_114;
wire n_0_115;
wire n_0_116;
wire n_0_117;
wire n_0_118;
wire n_0_119;
wire n_0_120;
wire opt_ipo_n23804;
wire slo__sro_n33778;
wire n_0_124;
wire n_0_0_2;
wire n_0_0_3;
wire n_0_0_4;
wire n_0_0_5;
wire n_0_0_6;
wire n_0_0_7;
wire n_0_0_8;
wire n_0_0_9;
wire n_0_0_10;
wire n_0_0_11;
wire n_0_0_12;
wire n_0_0_13;
wire n_0_0_14;
wire n_0_0_15;
wire n_0_0_16;
wire n_0_0_17;
wire n_0_0_18;
wire n_0_0_19;
wire n_0_0_20;
wire n_0_0_21;
wire n_0_0_22;
wire n_0_0_23;
wire n_0_0_24;
wire n_0_0_25;
wire n_0_0_26;
wire CLOCK_sgo__n47093;
wire n_0_0_28;
wire uc_0;
wire uc_1;
wire uc_2;
wire uc_3;
wire uc_4;
wire uc_5;
wire uc_6;
wire uc_7;
wire uc_8;
wire uc_9;
wire uc_10;
wire uc_11;
wire uc_12;
wire uc_13;
wire uc_14;
wire uc_15;
wire uc_16;
wire uc_17;
wire uc_18;
wire uc_19;
wire uc_20;
wire uc_21;
wire uc_22;
wire uc_23;
wire uc_24;
wire uc_25;
wire uc_26;
wire uc_27;
wire uc_28;
wire uc_29;
wire uc_30;
wire uc_31;
wire uc_32;
wire uc_33;
wire uc_34;
wire uc_35;
wire uc_36;
wire uc_37;
wire uc_38;
wire uc_39;
wire uc_40;
wire uc_41;
wire uc_42;
wire uc_43;
wire uc_44;
wire uc_45;
wire uc_46;
wire uc_47;
wire uc_48;
wire uc_49;
wire uc_50;
wire uc_51;
wire uc_52;
wire uc_53;
wire uc_54;
wire uc_55;
wire uc_56;
wire uc_57;
wire uc_58;
wire uc_59;
wire uc_60;
wire n_0;
wire n_1;
wire n_2;
wire n_3;
wire n_4;
wire n_5;
wire n_6;
wire n_7;
wire n_8;
wire n_9;
wire n_10;
wire n_11;
wire n_12;
wire n_13;
wire n_14;
wire n_15;
wire n_16;
wire n_17;
wire n_18;
wire n_19;
wire n_20;
wire n_21;
wire n_22;
wire n_23;
wire n_24;
wire n_25;
wire n_26;
wire n_27;
wire n_28;
wire n_29;
wire n_30;
wire n_31;
wire n_32;
wire n_33;
wire n_34;
wire n_35;
wire n_36;
wire n_37;
wire n_38;
wire n_39;
wire n_40;
wire n_41;
wire n_42;
wire n_43;
wire n_44;
wire n_45;
wire n_46;
wire n_47;
wire n_48;
wire n_49;
wire n_50;
wire n_51;
wire n_52;
wire CLOCK_slo__n54661;
wire n_54;
wire n_55;
wire n_56;
wire n_57;
wire CLOCK_slo__sro_n50363;
wire CLOCK_slo__sro_n51620;
wire slo__sro_n33466;
wire slo__mro_n33299;
wire CLOCK_slo__sro_n62669;
wire uc_61;
wire uc_62;
wire hfn_ipo_n25;
wire hfn_ipo_n26;
wire hfn_ipo_n27;
wire slo__sro_n35198;
wire hfn_ipo_n29;
wire hfn_ipo_n30;
wire hfn_ipo_n31;
wire hfn_ipo_n32;
wire hfn_ipo_n33;
wire hfn_ipo_n34;
wire hfn_ipo_n35;
wire hfn_ipo_n36;
wire sgo__n1292;
wire sgo__n1314;
wire sgo__n1306;
wire sgo__sro_n1582;
wire sgo__n1271;
wire sgo__n1276;
wire sgo__n1311;
wire sgo__sro_n1583;
wire sgo__sro_n1584;
wire sgo__sro_n1599;
wire sgo__sro_n1600;
wire sgo__sro_n1601;
wire sgo__sro_n1213;
wire sgo__sro_n1214;
wire sgo__sro_n1215;
wire sgo__sro_n1644;
wire sgo__sro_n1645;
wire slo__n26761;
wire slo__n15087;
wire sgo__sro_n1676;
wire sgo__sro_n1557;
wire slo__n37415;
wire sgo__sro_n1559;
wire sgo__sro_n1686;
wire sgo__sro_n1687;
wire sgo__sro_n1688;
wire slo__sro_n2106;
wire slo__sro_n2107;
wire slo__sro_n2108;
wire slo__sro_n2123;
wire slo__sro_n2142;
wire slo__sro_n2143;
wire slo__sro_n2144;
wire slo__sro_n2164;
wire slo__sro_n2165;
wire slo__sro_n2166;
wire slo__sro_n2167;
wire slo__sro_n2195;
wire slo__sro_n2196;
wire slo__sro_n2207;
wire slo__sro_n2208;
wire slo__sro_n2209;
wire slo__sro_n2221;
wire slo__sro_n2222;
wire slo__sro_n2230;
wire slo__sro_n2231;
wire slo__sro_n2232;
wire slo__sro_n2243;
wire slo__sro_n2244;
wire slo__sro_n2252;
wire slo__sro_n2253;
wire slo__sro_n2260;
wire slo__sro_n2261;
wire slo__sro_n2262;
wire slo__sro_n2273;
wire slo__sro_n2274;
wire slo__sro_n2285;
wire slo__sro_n2286;
wire slo__sro_n2287;
wire slo__sro_n2307;
wire slo__sro_n2308;
wire slo__sro_n2309;
wire slo__sro_n2318;
wire slo__sro_n2319;
wire slo__sro_n2338;
wire slo__sro_n2339;
wire slo__sro_n2346;
wire slo__sro_n2347;
wire slo__sro_n2348;
wire slo__sro_n35271;
wire slo__sro_n2370;
wire slo__sro_n2371;
wire slo__sro_n2372;
wire slo__sro_n2401;
wire slo__sro_n2408;
wire slo__sro_n2409;
wire slo__sro_n2410;
wire slo__n2560;
wire slo__n2708;
wire slo__n37437;
wire slo__sro_n2968;
wire slo__sro_n2969;
wire slo__sro_n2970;
wire slo__sro_n3057;
wire slo__sro_n3058;
wire slo__sro_n3059;
wire slo__n3800;
wire slo__sro_n3749;
wire slo__sro_n3751;
wire slo__sro_n3750;
wire slo__n3796;
wire slo__n3804;
wire slo__n3834;
wire slo__sro_n3904;
wire slo__sro_n3860;
wire CLOCK_slo__sro_n61296;
wire slo__sro_n3862;
wire slo__sro_n4232;
wire slo__sro_n4233;
wire slo__sro_n4244;
wire slo__sro_n4245;
wire slo__sro_n4287;
wire slo__sro_n4288;
wire slo__sro_n4339;
wire slo__sro_n4340;
wire slo__sro_n4341;
wire slo__sro_n4530;
wire slo__sro_n4312;
wire slo__sro_n4313;
wire slo__sro_n4615;
wire slo__sro_n4616;
wire slo__n33292;
wire slo__sro_n4528;
wire slo__sro_n4618;
wire opt_ipo_n45132;
wire slo__sro_n4661;
wire slo__sro_n4673;
wire slo__sro_n4674;
wire slo__sro_n4750;
wire CLOCK_sgo__sro_n47135;
wire slo__sro_n4690;
wire slo__sro_n4691;
wire slo__sro_n4752;
wire slo__sro_n4775;
wire slo__sro_n4785;
wire slo__sro_n4786;
wire slo__sro_n4787;
wire slo__sro_n4815;
wire slo__sro_n4816;
wire slo__sro_n4844;
wire slo__sro_n4845;
wire slo__sro_n4846;
wire slo__sro_n4847;
wire slo__sro_n4881;
wire slo__sro_n4882;
wire slo__sro_n4883;
wire slo__sro_n4923;
wire slo__n4944;
wire CLOCK_slo__sro_n61786;
wire slo__sro_n5017;
wire sgo__n471;
wire slo__sro_n5027;
wire slo__n4958;
wire slo__sro_n5057;
wire slo__sro_n5058;
wire slo__sro_n5059;
wire sgo__n482;
wire slo__sro_n5075;
wire slo__sro_n5119;
wire slo__sro_n5120;
wire CLOCK_slo__sro_n61698;
wire slo__n16975;
wire slo__sro_n5225;
wire sgo__n495;
wire slo__sro_n5226;
wire slo__sro_n5227;
wire CLOCK_slo__mro_n63532;
wire slo__sro_n5270;
wire slo__sro_n5285;
wire slo__n5306;
wire sgo__n508;
wire slo__sro_n5332;
wire slo__sro_n5333;
wire CLOCK_slo__sro_n59844;
wire slo__sro_n5353;
wire slo__sro_n5354;
wire slo__sro_n5417;
wire sgo__n521;
wire sgo__n522;
wire slo___n5717;
wire slo__sro_n5630;
wire slo__sro_n5679;
wire slo__sro_n5712;
wire slo__sro_n5713;
wire CLOCK_slo__sro_n52005;
wire sgo__n535;
wire slo__sro_n5844;
wire slo__sro_n37210;
wire slo__sro_n5876;
wire slo__sro_n5794;
wire sgo__n544;
wire slo__sro_n5878;
wire slo__sro_n5908;
wire slo__sro_n5964;
wire slo__sro_n5945;
wire sgo__n553;
wire slo__sro_n5946;
wire slo__sro_n31654;
wire slo__sro_n5988;
wire slo__sro_n6021;
wire slo__sro_n6038;
wire slo__sro_n6039;
wire sgo__n566;
wire slo__sro_n6040;
wire slo__sro_n6041;
wire slo__sro_n6090;
wire slo__sro_n6161;
wire slo__sro_n6162;
wire sgo__n577;
wire slo__sro_n6163;
wire slo__sro_n6240;
wire slo__sro_n6191;
wire slo__sro_n6192;
wire slo__sro_n6193;
wire slo__sro_n6194;
wire slo__sro_n6242;
wire CLOCK_slo__sro_n64636;
wire sgo__n594;
wire slo__sro_n6366;
wire CLOCK_slo__n55073;
wire slo__sro_n6283;
wire slo__sro_n6368;
wire slo__sro_n6369;
wire slo__sro_n6370;
wire sgo__n607;
wire slo__sro_n6520;
wire sgo__n610;
wire slo__sro_n6521;
wire sgo__n613;
wire slo__sro_n6522;
wire slo__sro_n6503;
wire sgo__n618;
wire slo__sro_n6504;
wire sgo__n621;
wire slo__sro_n6505;
wire slo__sro_n6455;
wire slo__sro_n6456;
wire slo__sro_n6457;
wire sgo__n630;
wire slo__sro_n6506;
wire CLOCK_slo__sro_n60776;
wire slo__sro_n6577;
wire sgo__n637;
wire slo__sro_n6578;
wire slo__sro_n6579;
wire slo__sro_n40939;
wire sgo__n644;
wire sgo__n645;
wire slo__sro_n6636;
wire slo__sro_n6637;
wire slo__sro_n6638;
wire slo__sro_n6674;
wire slo__sro_n6675;
wire sgo__n656;
wire slo__sro_n6676;
wire sgo__n659;
wire slo__sro_n6690;
wire slo__sro_n6691;
wire slo___n7115;
wire sgo__n666;
wire slo__sro_n6707;
wire slo__sro_n6708;
wire slo__sro_n6790;
wire slo__sro_n6737;
wire sgo__n675;
wire sgo__n676;
wire slo__sro_n6817;
wire slo__sro_n6830;
wire slo__sro_n6762;
wire slo__sro_n6763;
wire slo__sro_n6764;
wire sgo__n687;
wire sgo__n688;
wire slo__sro_n6765;
wire sgo__n691;
wire slo__sro_n31799;
wire slo__sro_n6852;
wire slo__sro_n6871;
wire slo__sro_n6872;
wire slo__sro_n6899;
wire slo___n6965;
wire slo___n6972;
wire slo__sro_n7038;
wire slo__sro_n7098;
wire slo__sro_n7073;
wire sgo__n711;
wire slo__sro_n31655;
wire sgo__n714;
wire sgo__n715;
wire slo__sro_n7075;
wire slo__sro_n6955;
wire slo__sro_n7017;
wire slo__sro_n7018;
wire slo__sro_n7019;
wire slo__sro_n7020;
wire slo__sro_n7187;
wire slo__sro_n7188;
wire slo__sro_n7189;
wire slo__sro_n7309;
wire slo__sro_n7331;
wire slo__sro_n7332;
wire slo__sro_n7395;
wire slo__sro_n7407;
wire slo__sro_n7219;
wire CLOCK_sgo__sro_n47198;
wire slo__sro_n7333;
wire slo__sro_n7334;
wire slo__sro_n7408;
wire slo__sro_n7422;
wire slo__sro_n7436;
wire slo__sro_n7307;
wire slo__sro_n7308;
wire slo__sro_n7448;
wire slo__sro_n7465;
wire slo__sro_n7467;
wire slo__sro_n37482;
wire slo__sro_n7478;
wire slo__sro_n7633;
wire slo__sro_n7691;
wire slo__sro_n7708;
wire slo__n7753;
wire slo__sro_n7689;
wire slo__sro_n7515;
wire CLOCK_slo__sro_n49604;
wire slo__sro_n7773;
wire slo__sro_n7774;
wire slo__sro_n7557;
wire slo__sro_n7775;
wire slo__sro_n40937;
wire slo__sro_n7834;
wire slo__sro_n7835;
wire slo__sro_n7911;
wire slo__sro_n19450;
wire slo__sro_n7898;
wire slo__sro_n7899;
wire slo__sro_n7913;
wire CLOCK_sgo__sro_n47261;
wire slo__sro_n7933;
wire slo__sro_n7946;
wire slo__sro_n7947;
wire slo__sro_n7961;
wire CLOCK_slo__n53754;
wire slo__sro_n8028;
wire slo__sro_n8029;
wire slo__sro_n8030;
wire slo__sro_n8046;
wire slo__sro_n8047;
wire slo__sro_n8057;
wire slo__sro_n8092;
wire slo__sro_n8180;
wire drc_ipo_n26587;
wire slo__sro_n8245;
wire slo__sro_n8294;
wire slo__sro_n8295;
wire slo__sro_n8296;
wire slo__sro_n8297;
wire slo__sro_n8311;
wire slo___n8747;
wire slo__sro_n8338;
wire slo__sro_n8340;
wire slo__sro_n8356;
wire slo__sro_n8357;
wire slo__sro_n8358;
wire slo__sro_n8368;
wire slo__sro_n8369;
wire slo__sro_n8370;
wire slo__sro_n8380;
wire slo__sro_n8391;
wire slo__sro_n8392;
wire slo__sro_n8402;
wire slo__sro_n8403;
wire slo__sro_n8404;
wire slo__sro_n40007;
wire slo__sro_n8415;
wire slo__sro_n8416;
wire slo__sro_n8417;
wire slo__sro_n8431;
wire slo__sro_n8432;
wire slo__sro_n8450;
wire slo__sro_n8451;
wire slo__sro_n8452;
wire slo__sro_n8453;
wire slo__sro_n8581;
wire slo__sro_n8488;
wire slo__sro_n8489;
wire slo__sro_n8558;
wire slo__sro_n8559;
wire slo__sro_n8603;
wire slo__sro_n8604;
wire slo__sro_n8605;
wire slo__sro_n8669;
wire slo__sro_n8646;
wire slo__sro_n8685;
wire slo__sro_n8686;
wire CLOCK_slo__sro_n49672;
wire slo__sro_n8742;
wire slo__sro_n8776;
wire slo__sro_n8731;
wire slo__sro_n8764;
wire slo__sro_n8765;
wire slo__sro_n8766;
wire slo__sro_n8778;
wire slo__sro_n21436;
wire slo__sro_n8916;
wire slo__sro_n8917;
wire slo__sro_n8872;
wire slo__sro_n8873;
wire slo__sro_n8874;
wire slo__sro_n8875;
wire slo__sro_n8901;
wire slo__sro_n8902;
wire slo__sro_n8903;
wire slo__sro_n8919;
wire slo__sro_n8965;
wire slo__sro_n8949;
wire slo__sro_n8979;
wire slo__sro_n8992;
wire slo__sro_n8993;
wire slo__sro_n8994;
wire slo__sro_n9008;
wire slo__sro_n9009;
wire slo__sro_n9010;
wire slo__sro_n9029;
wire slo__sro_n9030;
wire slo__sro_n9086;
wire slo__sro_n9075;
wire slo__sro_n9123;
wire slo__sro_n9124;
wire slo__sro_n9165;
wire slo__sro_n9194;
wire slo__sro_n9195;
wire slo__sro_n9196;
wire slo__sro_n9197;
wire slo__sro_n9243;
wire slo__sro_n9244;
wire slo__sro_n9245;
wire CLOCK_sgo__sro_n47395;
wire slo__sro_n9429;
wire slo__sro_n22110;
wire slo__sro_n9390;
wire CLOCK_slo__sro_n48740;
wire slo__sro_n9469;
wire slo__sro_n9470;
wire slo__sro_n9471;
wire slo__sro_n9535;
wire slo__n27411;
wire slo__sro_n9672;
wire slo__sro_n9673;
wire slo__sro_n9711;
wire slo__sro_n20323;
wire slo__sro_n9753;
wire slo__sro_n9713;
wire slo__sro_n9805;
wire slo__sro_n9754;
wire slo__sro_n9755;
wire slo__sro_n9745;
wire slo__sro_n9756;
wire CLOCK_slo__sro_n51474;
wire CLOCK_slo__sro_n51387;
wire CLOCK_slo__sro_n51388;
wire slo__sro_n9794;
wire slo__sro_n9916;
wire slo__sro_n9873;
wire slo__sro_n9874;
wire slo__sro_n9875;
wire slo__sro_n9977;
wire slo__sro_n9978;
wire slo__sro_n9979;
wire CLOCK_sgo__sro_n47212;
wire slo__sro_n29380;
wire slo__sro_n27838;
wire slo__sro_n10080;
wire slo__sro_n10099;
wire slo__sro_n10100;
wire slo__n10168;
wire slo__sro_n34087;
wire CLOCK_slo__mro_n51371;
wire slo__sro_n10273;
wire slo__n10331;
wire slo__sro_n10379;
wire slo__sro_n10311;
wire slo__sro_n10650;
wire slo__sro_n10426;
wire slo__sro_n10428;
wire slo__sro_n10429;
wire slo__sro_n10370;
wire slo__sro_n34361;
wire slo__sro_n10560;
wire slo__sro_n10518;
wire slo__sro_n10561;
wire slo__sro_n10562;
wire slo__sro_n32470;
wire slo__sro_n10651;
wire slo__sro_n10652;
wire CLOCK_slo__sro_n60679;
wire slo__sro_n10674;
wire slo__n10634;
wire slo__sro_n10675;
wire slo__sro_n10676;
wire slo__sro_n10694;
wire slo__sro_n10713;
wire slo__n10734;
wire slo__sro_n10771;
wire slo__sro_n10772;
wire slo__sro_n11080;
wire CLOCK_slo__sro_n49662;
wire slo__sro_n10839;
wire slo__sro_n11124;
wire slo__sro_n11125;
wire slo__sro_n10956;
wire CLOCK_slo__sro_n50083;
wire slo__sro_n10905;
wire slo__n10929;
wire CLOCK_sgo__sro_n47761;
wire slo__sro_n11126;
wire slo__sro_n11034;
wire slo__sro_n11035;
wire slo__sro_n11071;
wire slo__n38018;
wire slo__sro_n11215;
wire slo__sro_n11216;
wire slo__mro_n33239;
wire slo__sro_n11218;
wire slo__n11164;
wire slo__sro_n11317;
wire slo__n11270;
wire slo__sro_n11318;
wire slo__sro_n11319;
wire slo__sro_n11383;
wire slo__n11427;
wire slo__sro_n11437;
wire slo__sro_n11438;
wire slo__sro_n11483;
wire slo__sro_n11473;
wire slo__sro_n37401;
wire slo__n11253;
wire slo__n11487;
wire slo__sro_n11496;
wire slo__sro_n11706;
wire slo__sro_n11596;
wire slo__sro_n11597;
wire slo__sro_n11707;
wire slo__n11671;
wire slo__n12473;
wire slo__sro_n11708;
wire slo__sro_n11633;
wire slo__sro_n11709;
wire slo__sro_n11728;
wire slo__sro_n11729;
wire slo__sro_n11755;
wire slo__sro_n11797;
wire slo__sro_n11798;
wire slo__sro_n11784;
wire slo__sro_n11785;
wire slo__sro_n11786;
wire slo__sro_n11799;
wire slo__sro_n11828;
wire slo__sro_n11829;
wire slo__sro_n11830;
wire slo__sro_n11831;
wire slo__sro_n42332;
wire slo__sro_n11872;
wire slo__n11990;
wire opt_ipo_n45121;
wire slo__n12005;
wire CLOCK_sgo__sro_n48086;
wire slo__sro_n11889;
wire slo__sro_n12060;
wire slo__n12071;
wire slo__sro_n12111;
wire slo__sro_n12112;
wire slo__sro_n12113;
wire slo__sro_n12224;
wire slo__n11938;
wire slo__n12190;
wire slo__n29395;
wire slo__sro_n12329;
wire slo__sro_n12226;
wire slo__sro_n12227;
wire slo__sro_n12255;
wire slo__sro_n12256;
wire slo__sro_n12257;
wire slo___n12846;
wire slo__sro_n12465;
wire slo__sro_n12491;
wire slo__sro_n12492;
wire slo__sro_n12493;
wire slo__sro_n12507;
wire slo__sro_n12508;
wire slo__sro_n12534;
wire slo__sro_n12524;
wire slo__sro_n12525;
wire slo__sro_n12557;
wire slo__sro_n12558;
wire slo__sro_n12568;
wire slo__sro_n12569;
wire slo__sro_n12570;
wire slo__sro_n12571;
wire slo__n12811;
wire slo__n12606;
wire slo__sro_n12743;
wire slo__sro_n12744;
wire slo__sro_n12745;
wire slo__sro_n12746;
wire slo__n12843;
wire slo__sro_n12865;
wire slo__n12943;
wire slo__sro_n12923;
wire slo__sro_n12924;
wire slo__sro_n12925;
wire slo__sro_n12926;
wire slo__n13053;
wire slo__sro_n22024;
wire slo__sro_n12963;
wire slo__sro_n15043;
wire slo___n13169;
wire slo__sro_n13278;
wire slo__sro_n13701;
wire slo__n13153;
wire slo___n13213;
wire slo__sro_n13232;
wire slo__sro_n13235;
wire slo__sro_n13233;
wire slo__sro_n13234;
wire slo__sro_n13332;
wire slo__n13303;
wire slo__sro_n13333;
wire slo__sro_n13318;
wire slo__sro_n13334;
wire slo__sro_n13335;
wire slo__sro_n13356;
wire slo__sro_n13357;
wire slo__sro_n13371;
wire slo__sro_n13372;
wire slo__sro_n13382;
wire slo__sro_n13383;
wire slo__sro_n13384;
wire slo__sro_n13385;
wire slo__sro_n13471;
wire slo__sro_n13472;
wire slo__n13417;
wire slo__sro_n13461;
wire slo__sro_n13474;
wire slo__n13438;
wire slo__sro_n13522;
wire slo__n13528;
wire CLOCK_slo__sro_n49244;
wire slo__sro_n13545;
wire slo__n13621;
wire slo__sro_n13700;
wire slo__n13501;
wire slo__n13570;
wire slo__n13610;
wire slo__sro_n13702;
wire slo__sro_n13703;
wire CLOCK_slo__sro_n52594;
wire slo__sro_n13738;
wire slo__n13728;
wire CLOCK_slo__sro_n60125;
wire slo__sro_n13740;
wire slo__n13851;
wire slo__n13838;
wire slo__n13910;
wire CLOCK_slo__sro_n60275;
wire slo__n13799;
wire slo___n13777;
wire CLOCK_slo__sro_n62131;
wire slo__n13864;
wire slo__n13903;
wire slo__sro_n13953;
wire slo__sro_n13954;
wire slo__sro_n13955;
wire slo__n14026;
wire slo__sro_n14083;
wire slo__n13933;
wire slo__n14019;
wire slo__n14037;
wire slo__sro_n21634;
wire slo__sro_n14082;
wire slo__sro_n14084;
wire slo__n14095;
wire slo__sro_n14163;
wire slo__n14104;
wire slo__n14113;
wire slo__n14126;
wire slo__sro_n14164;
wire slo__sro_n14165;
wire slo__n14143;
wire slo__sro_n14166;
wire slo__n14207;
wire slo__sro_n30704;
wire slo__sro_n35616;
wire slo__sro_n14275;
wire CLOCK_slo__sro_n65089;
wire slo__n14340;
wire slo__n14465;
wire slo__n39286;
wire slo__sro_n14501;
wire slo__sro_n14441;
wire slo__n14568;
wire slo__sro_n14522;
wire slo__sro_n14523;
wire slo__sro_n14524;
wire slo__sro_n14525;
wire slo__n14633;
wire slo__n14640;
wire slo__n14647;
wire slo__n14626;
wire slo__n14684;
wire slo__n14691;
wire slo__n39417;
wire CLOCK_opt_ipo_n45730;
wire slo__sro_n14742;
wire slo__n14709;
wire slo__n14766;
wire slo__sro_n14855;
wire slo__sro_n14856;
wire CLOCK_slo__sro_n54706;
wire slo__n14894;
wire CLOCK_slo__sro_n62843;
wire slo__sro_n14915;
wire slo__n14949;
wire slo___n15030;
wire slo___n15116;
wire slo__sro_n14967;
wire slo___n15411;
wire slo__sro_n15079;
wire slo__sro_n15109;
wire slo__sro_n15110;
wire slo__n15162;
wire slo__sro_n15183;
wire slo__sro_n15184;
wire slo__sro_n22415;
wire slo__sro_n15143;
wire slo__sro_n15144;
wire slo__sro_n15145;
wire slo__sro_n15200;
wire slo__n15246;
wire slo__sro_n15534;
wire slo__sro_n15342;
wire slo__n15271;
wire slo__sro_n15343;
wire slo__sro_n15380;
wire slo__sro_n15381;
wire slo__sro_n15382;
wire slo__n15241;
wire slo__n15420;
wire slo__n15443;
wire slo__sro_n15470;
wire slo__sro_n15471;
wire slo__sro_n15472;
wire slo__sro_n15482;
wire slo__sro_n15483;
wire slo__sro_n15484;
wire slo__sro_n15485;
wire slo__sro_n15587;
wire slo__sro_n15671;
wire slo__sro_n15685;
wire slo___n15724;
wire slo__sro_n15669;
wire slo__n26713;
wire slo__sro_n15686;
wire slo__sro_n15687;
wire slo__sro_n15701;
wire slo__sro_n15702;
wire slo__sro_n15703;
wire slo__sro_n21498;
wire slo__sro_n15779;
wire slo__sro_n15796;
wire slo___n16283;
wire slo__n15821;
wire slo__sro_n15831;
wire slo__n15745;
wire slo__sro_n15832;
wire slo__sro_n15955;
wire slo__n15903;
wire slo__n15879;
wire slo__sro_n15956;
wire slo__n15870;
wire slo__n16022;
wire slo__n15894;
wire slo__n15976;
wire slo__n15969;
wire slo__n16063;
wire slo__n16143;
wire slo__n15930;
wire CLOCK_slo__sro_n51473;
wire slo__sro_n16001;
wire slo__sro_n16002;
wire slo__sro_n16003;
wire slo__sro_n16215;
wire slo__sro_n16180;
wire slo__n16152;
wire slo__sro_n16181;
wire slo__sro_n16182;
wire slo__sro_n29823;
wire slo__sro_n16183;
wire slo__sro_n16217;
wire slo__sro_n16218;
wire slo__sro_n16242;
wire slo___n16308;
wire slo__n16267;
wire slo__n16280;
wire slo___n16361;
wire slo__n16348;
wire slo__n16450;
wire slo__n16392;
wire CLOCK_slo__sro_n50974;
wire slo__n16343;
wire slo__sro_n16886;
wire slo__n16524;
wire slo__n16550;
wire slo__n16529;
wire slo__n16413;
wire slo__n16608;
wire slo__n16557;
wire slo__n16796;
wire slo__n16747;
wire slo__n16572;
wire slo__n16706;
wire slo__n16791;
wire slo__n17041;
wire slo__n16774;
wire slo__n16984;
wire slo__n16871;
wire slo__n16864;
wire slo__sro_n16910;
wire slo__sro_n17056;
wire slo__n17020;
wire slo__sro_n17057;
wire slo__sro_n17058;
wire slo__n17088;
wire slo__sro_n17074;
wire slo__sro_n17075;
wire slo__sro_n17076;
wire slo__n17214;
wire slo__sro_n17254;
wire slo__sro_n17238;
wire slo__sro_n17255;
wire slo__sro_n17256;
wire slo__sro_n17239;
wire slo__sro_n17240;
wire slo__sro_n17241;
wire slo__n17290;
wire slo___n17582;
wire slo__sro_n17353;
wire slo__sro_n17330;
wire slo__n17378;
wire slo___n17633;
wire slo___n17474;
wire CLOCK_slo__sro_n59232;
wire slo__sro_n17598;
wire slo__n17399;
wire slo__n17416;
wire slo__n17575;
wire slo__sro_n17647;
wire slo__sro_n17646;
wire slo__n17619;
wire slo__sro_n17648;
wire slo__sro_n17649;
wire slo__n17671;
wire slo__sro_n17782;
wire slo__n17680;
wire slo__sro_n17693;
wire slo__n17737;
wire slo__n17744;
wire slo__sro_n17761;
wire slo___n17886;
wire slo__sro_n17781;
wire slo__sro_n18042;
wire slo__n17821;
wire slo__sro_n17951;
wire slo__n17921;
wire CLOCK_slo__sro_n51512;
wire slo__sro_n17953;
wire slo___n18137;
wire slo__n17942;
wire slo__n18019;
wire slo__n18084;
wire slo__sro_n18043;
wire slo__sro_n18044;
wire slo__sro_n18343;
wire spw__n69100;
wire slo__n18297;
wire slo__sro_n18154;
wire slo__n18122;
wire slo__sro_n18155;
wire slo__sro_n18156;
wire slo__n18178;
wire slo__n18277;
wire CLOCK_slo__sro_n57702;
wire slo__n18653;
wire slo__n18328;
wire slo__sro_n18404;
wire slo__sro_n18405;
wire slo__sro_n18406;
wire slo__sro_n18480;
wire slo__sro_n18481;
wire CLOCK_slo__sro_n64638;
wire slo__sro_n18492;
wire slo__n18727;
wire slo__n18523;
wire slo___n18581;
wire slo__n18732;
wire slo__n18626;
wire slo__n18737;
wire CLOCK_sgo__sro_n47338;
wire slo__n18771;
wire slo__n18766;
wire slo__n18776;
wire slo__n18930;
wire slo__sro_n18863;
wire slo__sro_n18951;
wire slo__n18942;
wire slo__n18848;
wire slo__n18877;
wire slo___n19273;
wire slo__n19067;
wire slo__n18973;
wire slo__n18982;
wire slo__n18991;
wire slo__sro_n19076;
wire slo__sro_n19077;
wire slo__sro_n19078;
wire slo__sro_n19024;
wire slo__sro_n19025;
wire slo__sro_n19026;
wire slo__sro_n19027;
wire slo___n19182;
wire slo__n19102;
wire slo__sro_n19349;
wire slo__n19282;
wire slo__sro_n19351;
wire slo__n19179;
wire slo__sro_n19383;
wire slo__n19255;
wire slo__sro_n19350;
wire slo__n19320;
wire slo__sro_n19384;
wire slo__sro_n19385;
wire slo__sro_n19420;
wire slo__sro_n19421;
wire slo__sro_n19422;
wire slo__sro_n19423;
wire slo__sro_n19437;
wire slo__sro_n19438;
wire slo__sro_n19439;
wire slo__sro_n19567;
wire slo__sro_n19543;
wire slo__sro_n19544;
wire slo__sro_n19545;
wire slo__sro_n19546;
wire slo__sro_n19569;
wire slo__sro_n19570;
wire slo__sro_n19727;
wire slo__sro_n19728;
wire slo__sro_n19839;
wire slo__sro_n19627;
wire slo__sro_n19628;
wire slo__sro_n19753;
wire slo__sro_n19754;
wire slo__sro_n19971;
wire slo__sro_n19751;
wire slo__sro_n19807;
wire slo__sro_n19808;
wire slo__sro_n19972;
wire slo__sro_n19673;
wire slo__sro_n19674;
wire slo__sro_n19675;
wire slo__sro_n19676;
wire slo__sro_n19958;
wire slo__sro_n19959;
wire slo__sro_n19894;
wire slo__sro_n19895;
wire slo__sro_n19896;
wire slo__sro_n19897;
wire slo__sro_n19998;
wire slo__sro_n19999;
wire slo__sro_n20000;
wire slo__sro_n20067;
wire slo__sro_n20068;
wire CLOCK_slo__n60586;
wire slo__sro_n20056;
wire slo__sro_n20057;
wire slo__sro_n20058;
wire slo__sro_n20081;
wire slo__sro_n20146;
wire slo__sro_n20147;
wire slo__sro_n20261;
wire slo__sro_n20262;
wire slo__sro_n32484;
wire slo__sro_n20127;
wire slo__sro_n20285;
wire slo__sro_n20286;
wire slo__sro_n20287;
wire slo__sro_n20288;
wire slo__sro_n20324;
wire slo__sro_n20395;
wire slo__sro_n20396;
wire slo__sro_n20420;
wire slo__sro_n20506;
wire slo__mro_n33267;
wire slo__mro_n33266;
wire slo__sro_n20472;
wire slo__sro_n20473;
wire slo__sro_n20474;
wire slo__sro_n20475;
wire CLOCK_sgo__sro_n47394;
wire CLOCK_sgo__sro_n47199;
wire slo__sro_n20568;
wire slo__sro_n20614;
wire slo__sro_n20615;
wire slo__sro_n20680;
wire slo__sro_n20681;
wire slo__sro_n20682;
wire slo__sro_n20683;
wire slo__sro_n20735;
wire slo__sro_n20817;
wire slo__sro_n20818;
wire slo__sro_n20819;
wire slo__sro_n20820;
wire slo__sro_n20846;
wire slo__sro_n20847;
wire slo__sro_n20848;
wire slo__sro_n20886;
wire slo__sro_n20887;
wire slo__sro_n20888;
wire slo__sro_n20913;
wire slo__sro_n20914;
wire slo__sro_n20915;
wire slo__sro_n20924;
wire slo__sro_n21011;
wire slo__sro_n21012;
wire slo__sro_n21212;
wire slo__sro_n21314;
wire slo__sro_n21315;
wire slo__sro_n21316;
wire slo__sro_n21317;
wire CLOCK_slo__sro_n62825;
wire slo__sro_n20974;
wire slo__sro_n21346;
wire slo__sro_n21347;
wire slo__sro_n21348;
wire slo__sro_n21349;
wire slo__sro_n21380;
wire slo__sro_n21381;
wire slo__sro_n21382;
wire slo__sro_n21438;
wire slo__sro_n21439;
wire slo__sro_n21499;
wire slo__sro_n21500;
wire slo__sro_n21560;
wire slo__sro_n21561;
wire slo__sro_n21633;
wire slo__sro_n40960;
wire slo__sro_n21603;
wire slo__sro_n21635;
wire slo__sro_n21663;
wire slo__sro_n21664;
wire slo__sro_n21665;
wire CLOCK_slo___n64354;
wire slo__sro_n21678;
wire slo__sro_n21753;
wire slo__sro_n21754;
wire slo__sro_n21755;
wire drc_ipo_n26586;
wire slo__sro_n21796;
wire slo__sro_n21797;
wire slo__sro_n21836;
wire slo__sro_n21941;
wire slo__sro_n21940;
wire slo__sro_n21942;
wire slo__sro_n22025;
wire slo__sro_n22026;
wire slo__sro_n22111;
wire slo__sro_n22112;
wire slo__sro_n22113;
wire slo__sro_n22133;
wire slo__sro_n22134;
wire slo__sro_n22326;
wire slo__sro_n22327;
wire slo__sro_n22328;
wire slo__mro_n33031;
wire slo__mro_n33030;
wire slo__sro_n22350;
wire slo__sro_n22416;
wire slo__sro_n22417;
wire slo__sro_n22432;
wire slo__sro_n22433;
wire slo__sro_n22458;
wire CLOCK_slo__sro_n62512;
wire CLOCK_slo__sro_n62513;
wire slo__sro_n22580;
wire slo__sro_n22553;
wire slo__sro_n22554;
wire slo__sro_n22555;
wire slo__sro_n22624;
wire slo__sro_n22625;
wire slo__sro_n22701;
wire slo__sro_n22677;
wire slo__sro_n22678;
wire slo__sro_n22679;
wire slo__sro_n22703;
wire slo__sro_n22736;
wire slo__sro_n22743;
wire slo__sro_n22744;
wire slo__sro_n22745;
wire slo__sro_n22779;
wire slo__sro_n22769;
wire slo__sro_n22770;
wire slo__sro_n22771;
wire slo__sro_n22780;
wire slo__sro_n22781;
wire slo__sro_n22782;
wire slo__sro_n22874;
wire slo__sro_n22875;
wire slo__sro_n22964;
wire slo__sro_n22965;
wire slo__sro_n23158;
wire CLOCK_slo__n53479;
wire slo__sro_n23125;
wire slo__sro_n23160;
wire slo___n23218;
wire slo___n23221;
wire slo___n23226;
wire slo___n23229;
wire slo___n23232;
wire slo___n23235;
wire drc_ipo_n26573;
wire slo___n23239;
wire slo___n23244;
wire slo___n23247;
wire slo___n23268;
wire drc_ipo_n26577;
wire slo___n23274;
wire slo___n23277;
wire drc_ipo_n26574;
wire slo___n23353;
wire slo__n23262;
wire slo__n23263;
wire spt__n66415;
wire slo___n23359;
wire slo___n23364;
wire slo___n23367;
wire slo___n23404;
wire slo___n23407;
wire slo___n23430;
wire slo__n23298;
wire slo__n23299;
wire slo___n23451;
wire drc_ipo_n26575;
wire slo___n23457;
wire CLOCK_slo__sro_n61284;
wire slo___n23463;
wire slo___n23466;
wire slo__n23424;
wire slo__n23425;
wire slo__n23445;
wire slo__n23446;
wire drc_ipo_n26609;
wire slo__n23398;
wire slo__n23399;
wire drc_ipo_n26610;
wire CLOCK_sgo__n46808;
wire drc_ipo_n26613;
wire drc_ipo_n26614;
wire drc_ipo_n26615;
wire drc_ipo_n26616;
wire drc_ipo_n26617;
wire drc_ipo_n26618;
wire drc_ipo_n26620;
wire drc_ipo_n26621;
wire drc_ipo_n26624;
wire drc_ipo_n26625;
wire CLOCK_slo__sro_n62842;
wire CLOCK_slo__sro_n62786;
wire slo__n26638;
wire CLOCK_slo__sro_n62785;
wire CLOCK_slo__sro_n62784;
wire spt__n66349;
wire CLOCK_slo__sro_n62746;
wire CLOCK_slo__sro_n62745;
wire CLOCK_slo__sro_n62783;
wire slo__n26645;
wire opt_ipo_n23872;
wire slo__n28104;
wire slo__n26648;
wire CLOCK_slo__sro_n62530;
wire CLOCK_slo__mro_n62208;
wire CLOCK_slo__sro_n62129;
wire CLOCK_slo__sro_n61963;
wire CLOCK_slo__sro_n61962;
wire slo__n26654;
wire CLOCK_slo__sro_n61944;
wire CLOCK_slo__sro_n61396;
wire CLOCK_slo__sro_n61945;
wire slo__n26658;
wire CLOCK_slo__sro_n61943;
wire CLOCK_sgo__n47094;
wire slo__n26805;
wire slo__sro_n27140;
wire slo__sro_n27583;
wire slo__sro_n26911;
wire slo__sro_n27159;
wire slo__sro_n27251;
wire slo__sro_n27252;
wire slo__n27410;
wire slo__sro_n27160;
wire slo__sro_n27392;
wire slo__n26894;
wire slo__n26895;
wire slo__n26896;
wire slo__sro_n27138;
wire slo__sro_n27253;
wire slo__sro_n27360;
wire slo__sro_n27361;
wire slo__sro_n27362;
wire slo__sro_n27499;
wire slo__sro_n27500;
wire slo__sro_n27501;
wire slo__sro_n27339;
wire slo__sro_n27571;
wire slo__sro_n27572;
wire slo__sro_n27573;
wire slo__sro_n27584;
wire slo__sro_n27691;
wire CLOCK_sgo__sro_n47211;
wire CLOCK_slo__mro_n63339;
wire slo__sro_n27726;
wire slo__sro_n27728;
wire slo__sro_n27862;
wire slo__sro_n27690;
wire slo__sro_n27972;
wire slo__sro_n27891;
wire slo__sro_n27892;
wire slo__sro_n27893;
wire slo__sro_n27973;
wire slo__sro_n27822;
wire slo__sro_n27823;
wire slo__sro_n27974;
wire slo__sro_n28007;
wire slo__sro_n28008;
wire slo__n28070;
wire slo__n28071;
wire slo__n28105;
wire slo__sro_n28181;
wire slo__sro_n28182;
wire slo__sro_n28183;
wire slo__sro_n28285;
wire slo__sro_n28421;
wire slo__sro_n28524;
wire slo__sro_n28333;
wire slo__sro_n28334;
wire slo__sro_n28525;
wire slo__sro_n28526;
wire slo__sro_n28564;
wire slo__sro_n28422;
wire slo__sro_n28283;
wire slo__sro_n28284;
wire slo__n28539;
wire opt_ipo_n24063;
wire slo__sro_n29018;
wire slo__sro_n29019;
wire slo__sro_n28659;
wire slo__sro_n28660;
wire opt_ipo_n24075;
wire slo__sro_n28775;
wire slo__sro_n28989;
wire slo__sro_n28776;
wire slo__sro_n28990;
wire slo__sro_n29068;
wire slo__sro_n29069;
wire slo__sro_n28777;
wire slo__sro_n29225;
wire slo__sro_n29226;
wire slo__sro_n29176;
wire slo__sro_n29228;
wire slo__sro_n29365;
wire slo__sro_n29205;
wire slo__sro_n29206;
wire slo__sro_n29207;
wire slo__sro_n29227;
wire slo__sro_n29363;
wire slo__sro_n29381;
wire slo__sro_n29444;
wire slo__sro_n29693;
wire slo__sro_n29651;
wire slo__sro_n29675;
wire slo__sro_n29650;
wire slo__sro_n29489;
wire slo__sro_n29490;
wire slo__sro_n29491;
wire slo__sro_n29676;
wire slo__sro_n29677;
wire slo__sro_n29523;
wire slo__sro_n29524;
wire slo__sro_n29525;
wire slo__sro_n29526;
wire slo__sro_n30018;
wire slo__sro_n29822;
wire CLOCK_sgo__sro_n47245;
wire slo__sro_n29773;
wire opt_ipo_n45107;
wire opt_ipo_n24166;
wire slo__sro_n29824;
wire slo__sro_n29858;
wire CLOCK_slo__sro_n64639;
wire opt_ipo_n24173;
wire slo__sro_n29860;
wire slo__sro_n29881;
wire CLOCK_sgo__sro_n47134;
wire slo__sro_n29917;
wire slo__sro_n29918;
wire slo__sro_n29919;
wire opt_ipo_n24190;
wire slo__sro_n30020;
wire slo__sro_n30033;
wire opt_ipo_n24196;
wire slo__sro_n30034;
wire slo__sro_n30284;
wire slo__sro_n30110;
wire slo__sro_n30111;
wire slo__sro_n30145;
wire slo__sro_n30071;
wire slo__sro_n30072;
wire slo__sro_n30073;
wire slo__sro_n30112;
wire slo__sro_n30113;
wire slo__sro_n30147;
wire slo__sro_n30286;
wire slo__sro_n30207;
wire slo__sro_n30208;
wire slo__sro_n30209;
wire slo__sro_n30264;
wire slo__sro_n30265;
wire slo__sro_n30266;
wire slo__sro_n30287;
wire slo__n30589;
wire slo__n30670;
wire slo__sro_n30362;
wire opt_ipo_n24251;
wire slo__sro_n30364;
wire slo__sro_n31362;
wire slo__sro_n30504;
wire slo__sro_n30505;
wire slo__sro_n30506;
wire slo__sro_n31363;
wire slo__sro_n37221;
wire slo__sro_n30706;
wire CLOCK_sgo__sro_n47150;
wire slo__sro_n30996;
wire slo__sro_n30921;
wire slo__sro_n30922;
wire slo__sro_n30923;
wire slo__sro_n30924;
wire opt_ipo_n24285;
wire slo__sro_n30998;
wire slo__sro_n31053;
wire slo__sro_n31088;
wire slo__sro_n31089;
wire slo__sro_n31220;
wire slo__sro_n31218;
wire slo__sro_n31234;
wire slo__sro_n31235;
wire slo__sro_n31236;
wire slo__sro_n31237;
wire slo__sro_n31559;
wire slo__sro_n31306;
wire slo__sro_n31307;
wire CLOCK_opt_ipo_n45742;
wire slo__mro_n31601;
wire slo__sro_n31560;
wire slo__sro_n31483;
wire opt_ipo_n24326;
wire slo__sro_n31484;
wire CLOCK_sgo__sro_n47148;
wire slo__sro_n31561;
wire slo__sro_n31562;
wire slo__sro_n31644;
wire slo__sro_n31645;
wire slo__sro_n31646;
wire slo__sro_n31657;
wire slo__sro_n31671;
wire slo__sro_n31672;
wire slo__n31700;
wire slo__sro_n31816;
wire opt_ipo_n24358;
wire slo__sro_n31800;
wire slo__sro_n31801;
wire slo__sro_n31818;
wire slo__sro_n31819;
wire slo__sro_n31831;
wire slo__sro_n31832;
wire slo__sro_n32028;
wire slo__sro_n32029;
wire slo__sro_n32026;
wire slo__sro_n32045;
wire slo__sro_n32046;
wire CLOCK_sgo__sro_n47197;
wire slo__sro_n32118;
wire slo__sro_n32119;
wire slo__sro_n32120;
wire CLOCK_slo__sro_n62931;
wire slo__sro_n32140;
wire slo__sro_n32182;
wire slo__sro_n32163;
wire slo__sro_n32164;
wire slo__sro_n32165;
wire slo__sro_n32166;
wire slo__sro_n32183;
wire slo__sro_n32184;
wire slo__sro_n32185;
wire slo__sro_n32204;
wire slo__sro_n32213;
wire slo__sro_n32316;
wire opt_ipo_n24431;
wire slo__sro_n32318;
wire opt_ipo_n45138;
wire slo__sro_n32357;
wire slo__sro_n32358;
wire slo__n32451;
wire slo__sro_n38698;
wire slo__sro_n32472;
wire slo__sro_n32473;
wire slo__sro_n32716;
wire slo__sro_n32717;
wire slo__mro_n33269;
wire slo__mro_n33268;
wire slo__mro_n33301;
wire slo__mro_n33302;
wire slo__sro_n33598;
wire slo__sro_n33789;
wire slo__sro_n34622;
wire slo__sro_n33526;
wire slo__sro_n33373;
wire slo__sro_n33527;
wire slo__sro_n34034;
wire slo__sro_n34035;
wire slo__sro_n34608;
wire slo__sro_n34247;
wire slo__sro_n34248;
wire slo__sro_n33677;
wire slo__sro_n34609;
wire slo__sro_n34756;
wire opt_ipo_n24503;
wire slo__sro_n34623;
wire CLOCK_slo__sro_n51957;
wire slo__sro_n34758;
wire slo__sro_n34940;
wire slo__sro_n33384;
wire slo__mro_n33237;
wire CLOCK_slo__sro_n58764;
wire slo__sro_n35378;
wire slo__sro_n35466;
wire slo__sro_n35617;
wire slo__sro_n35312;
wire slo__sro_n35313;
wire slo__mro_n33238;
wire slo__mro_n33014;
wire opt_ipo_n24541;
wire slo__sro_n35249;
wire slo__sro_n35250;
wire slo__sro_n34941;
wire slo__sro_n35145;
wire slo__n35114;
wire slo__n35115;
wire CLOCK_sgo__sro_n47263;
wire slo__sro_n35375;
wire slo__sro_n35376;
wire slo__sro_n35377;
wire slo__sro_n35618;
wire CLOCK_slo__sro_n50432;
wire slo__sro_n35419;
wire slo__sro_n36418;
wire slo__sro_n28286;
wire slo__sro_n28523;
wire slo__sro_n36417;
wire slo__sro_n36479;
wire slo__sro_n34095;
wire slo__sro_n34607;
wire slo__sro_n34126;
wire slo__sro_n34317;
wire slo__sro_n34606;
wire spt__n66327;
wire CLOCK_slo__sro_n61394;
wire slo__sro_n36419;
wire slo__sro_n36837;
wire slo__sro_n35681;
wire slo__sro_n35682;
wire slo__sro_n35683;
wire slo__sro_n35684;
wire slo__sro_n36088;
wire slo__sro_n35199;
wire CLOCK_slo__n60839;
wire slo__sro_n36567;
wire slo__sro_n36946;
wire slo__sro_n37222;
wire slo__sro_n36684;
wire slo__sro_n37092;
wire slo__sro_n37211;
wire slo__sro_n36913;
wire slo__sro_n36836;
wire slo__n35732;
wire slo__sro_n36944;
wire slo__sro_n36810;
wire slo__sro_n36933;
wire slo__sro_n37306;
wire slo__sro_n37223;
wire slo__sro_n36260;
wire slo__n36214;
wire slo__sro_n37053;
wire slo__sro_n37054;
wire slo__sro_n37055;
wire slo__sro_n37224;
wire slo__sro_n37307;
wire slo__sro_n37308;
wire slo__sro_n37390;
wire slo__sro_n37402;
wire slo__sro_n37403;
wire slo__sro_n37387;
wire slo__sro_n37388;
wire slo__sro_n37404;
wire slo__sro_n37405;
wire CLOCK_slo__sro_n49773;
wire opt_ipo_n24698;
wire slo__sro_n37483;
wire slo__n37463;
wire slo__sro_n37452;
wire opt_ipo_n24707;
wire slo__sro_n37454;
wire slo__sro_n37484;
wire slo__sro_n37485;
wire slo__n37502;
wire slo__sro_n37540;
wire opt_ipo_n24721;
wire slo__sro_n37842;
wire opt_ipo_n24727;
wire slo__n37528;
wire slo__sro_n38411;
wire slo__n38056;
wire slo__sro_n37843;
wire slo__sro_n36308;
wire slo__sro_n37999;
wire opt_ipo_n24743;
wire slo__sro_n36045;
wire slo__sro_n38408;
wire slo__n38227;
wire slo__n38240;
wire slo__n38193;
wire slo__sro_n38409;
wire slo__sro_n38324;
wire slo__sro_n38745;
wire slo__n38599;
wire slo__sro_n38410;
wire slo__sro_n38298;
wire slo__sro_n38299;
wire slo__sro_n38300;
wire CLOCK_slo__sro_n50186;
wire slo__n38566;
wire opt_ipo_n24784;
wire slo__sro_n38684;
wire slo__sro_n38685;
wire slo__sro_n38686;
wire slo__sro_n38687;
wire slo__sro_n37841;
wire CLOCK_slo__sro_n49188;
wire slo__sro_n38746;
wire slo__sro_n38747;
wire slo__sro_n38759;
wire slo__sro_n38760;
wire slo__sro_n38761;
wire slo__n38783;
wire slo__sro_n38915;
wire slo__sro_n38941;
wire slo__sro_n38942;
wire slo__sro_n38916;
wire slo__sro_n38807;
wire slo__sro_n38808;
wire CLOCK_sgo__sro_n47200;
wire slo__n38840;
wire slo__n38973;
wire slo__sro_n38943;
wire slo__n39285;
wire slo__n39136;
wire slo__n39084;
wire slo__sro_n39249;
wire slo__n39345;
wire slo__sro_n39122;
wire slo__sro_n39872;
wire slo__n39719;
wire slo__sro_n39363;
wire opt_ipo_n24861;
wire slo__sro_n39888;
wire slo__sro_n39768;
wire slo__sro_n39597;
wire slo__sro_n39513;
wire slo__sro_n39769;
wire slo__sro_n39770;
wire slo__sro_n39797;
wire slo__sro_n39889;
wire slo__sro_n39900;
wire slo__n39745;
wire slo__sro_n40961;
wire slo__sro_n39898;
wire slo__sro_n40008;
wire slo__sro_n40009;
wire slo__sro_n40010;
wire slo__n39957;
wire CLOCK_slo__sro_n49712;
wire slo__sro_n40292;
wire slo__n40090;
wire slo__n40097;
wire slo___n43257;
wire slo__sro_n40936;
wire slo__sro_n41807;
wire slo__sro_n41833;
wire CLOCK_slo__sro_n55084;
wire slo__sro_n40148;
wire slo__sro_n40149;
wire slo__sro_n40150;
wire slo__sro_n40938;
wire slo__sro_n41808;
wire slo__sro_n41144;
wire slo__sro_n41030;
wire CLOCK_slo__n65456;
wire slo__sro_n40371;
wire slo__sro_n41031;
wire slo__sro_n41029;
wire slo__sro_n41060;
wire slo__sro_n40769;
wire slo__sro_n40459;
wire spw__n67799;
wire slo__sro_n40462;
wire opt_ipo_n24966;
wire slo__sro_n41478;
wire CLOCK_sgo__sro_n47337;
wire slo__sro_n41809;
wire slo__sro_n41830;
wire slo__n41747;
wire slo__sro_n41831;
wire slo__sro_n41832;
wire slo__sro_n41810;
wire slo___n43247;
wire slo__sro_n42331;
wire CLOCK_opt_ipo_n45803;
wire CLOCK_sgo__sro_n47339;
wire CLOCK_opt_ipo_n45807;
wire CLOCK_slo__sro_n61297;
wire opt_ipo_n25006;
wire opt_ipo_n25007;
wire CLOCK_sgo__n46814;
wire opt_ipo_n45134;
wire CLOCK_opt_ipo_n45779;
wire opt_ipo_n43935;
wire CLOCK_sgo__n46815;
wire CLOCK_opt_ipo_n45825;
wire spt__n66340;
wire CLOCK_sgo__sro_n47296;
wire opt_ipo_n45144;
wire opt_ipo_n45145;
wire slo___n43254;
wire CLOCK_slo__sro_n64581;
wire CLOCK_sgo__sro_n47307;
wire CLOCK_sgo__sro_n47468;
wire CLOCK_sgo__sro_n47440;
wire CLOCK_sgo__n46841;
wire CLOCK_sgo__sro_n47298;
wire CLOCK_slo__sro_n59282;
wire CLOCK_slo__sro_n62894;
wire CLOCK_sgo__sro_n47441;
wire CLOCK_sgo__sro_n47442;
wire CLOCK_sgo__sro_n47469;
wire CLOCK_sgo__sro_n47470;
wire CLOCK_sgo__sro_n47501;
wire CLOCK_sgo__sro_n47502;
wire CLOCK_sgo__sro_n47503;
wire CLOCK_sgo__sro_n47538;
wire CLOCK_sgo__sro_n47562;
wire CLOCK_sgo__sro_n47539;
wire CLOCK_sgo__sro_n47540;
wire CLOCK_sgo__sro_n47541;
wire CLOCK_sgo__sro_n47560;
wire CLOCK_opt_ipo_n45873;
wire CLOCK_sgo__sro_n47592;
wire CLOCK_sgo__sro_n47593;
wire CLOCK_sgo__sro_n47602;
wire CLOCK_sgo__sro_n47603;
wire CLOCK_sgo__sro_n47604;
wire CLOCK_sgo__sro_n47621;
wire CLOCK_sgo__sro_n47622;
wire CLOCK_sgo__sro_n47623;
wire CLOCK_opt_ipo_n45736;
wire opt_ipo_n25116;
wire CLOCK_opt_ipo_n45894;
wire opt_ipo_n25120;
wire CLOCK_sgo__sro_n47111;
wire CLOCK_sgo__sro_n47682;
wire CLOCK_sgo__sro_n47683;
wire CLOCK_sgo__sro_n47701;
wire CLOCK_opt_ipo_n45906;
wire CLOCK_sgo__sro_n47733;
wire CLOCK_sgo__sro_n47734;
wire CLOCK_sgo__n48008;
wire CLOCK_opt_ipo_n45918;
wire CLOCK_sgo__n48011;
wire CLOCK_sgo__sro_n47762;
wire CLOCK_sgo__sro_n47798;
wire CLOCK_sgo__sro_n47799;
wire CLOCK_sgo__sro_n47800;
wire opt_ipo_n44105;
wire CLOCK_sgo__sro_n47822;
wire CLOCK_sgo__n46922;
wire CLOCK_slo__sro_n61348;
wire CLOCK_sgo__sro_n47823;
wire opt_ipo_n44116;
wire CLOCK_sgo__sro_n47825;
wire CLOCK_sgo__sro_n47835;
wire CLOCK_sgo__sro_n47836;
wire CLOCK_sgo__n46934;
wire CLOCK_sgo__sro_n47837;
wire CLOCK_sgo__n46937;
wire CLOCK_sgo__sro_n47846;
wire CLOCK_sgo__sro_n47847;
wire CLOCK_sgo__n46942;
wire CLOCK_sgo__sro_n48087;
wire CLOCK_opt_ipo_n45969;
wire CLOCK_slo__sro_n48338;
wire CLOCK_slo__n48430;
wire CLOCK_sgo__n46950;
wire CLOCK_opt_ipo_n45978;
wire opt_ipo_n45366;
wire CLOCK_sgo__sro_n48189;
wire CLOCK_sgo__sro_n48190;
wire CLOCK_slo__sro_n62930;
wire CLOCK_slo__sro_n48636;
wire CLOCK_slo__sro_n64637;
wire CLOCK_slo__sro_n48699;
wire CLOCK_slo__sro_n48741;
wire CLOCK_slo__sro_n48742;
wire CLOCK_slo__sro_n48812;
wire CLOCK_slo__sro_n48814;
wire spw__n69101;
wire CLOCK_opt_ipo_n46005;
wire CLOCK_slo__sro_n48874;
wire CLOCK_slo__sro_n48784;
wire CLOCK_slo__sro_n48785;
wire CLOCK_slo__sro_n48786;
wire CLOCK_slo__sro_n48875;
wire CLOCK_slo__sro_n48876;
wire CLOCK_slo__n48906;
wire CLOCK_slo__sro_n48960;
wire CLOCK_slo__sro_n48976;
wire spw__n67656;
wire CLOCK_opt_ipo_n46029;
wire CLOCK_slo__sro_n48978;
wire CLOCK_slo__sro_n49022;
wire CLOCK_slo__sro_n49023;
wire CLOCK_opt_ipo_n46038;
wire CLOCK_sgo__n47002;
wire CLOCK_sgo__n47003;
wire CLOCK_sgo__n47004;
wire CLOCK_sgo__n47005;
wire CLOCK_slo__sro_n49024;
wire CLOCK_slo__sro_n49025;
wire CLOCK_slo__n49050;
wire CLOCK_slo__sro_n49084;
wire CLOCK_slo__sro_n49120;
wire CLOCK_slo__sro_n49121;
wire CLOCK_slo__n49140;
wire CLOCK_slo__n49141;
wire CLOCK_slo__sro_n62130;
wire CLOCK_slo__sro_n62128;
wire CLOCK_slo__sro_n62488;
wire CLOCK_sgo__n47025;
wire CLOCK_slo__sro_n61395;
wire opt_ipo_n45480;
wire CLOCK_slo__sro_n49189;
wire CLOCK_slo__sro_n49190;
wire CLOCK_slo__sro_n49191;
wire CLOCK_slo__sro_n49216;
wire CLOCK_slo__sro_n49217;
wire CLOCK_slo__sro_n49218;
wire CLOCK_slo__sro_n49069;
wire CLOCK_slo__sro_n49348;
wire CLOCK_slo__sro_n49349;
wire CLOCK_sgo__n47049;
wire CLOCK_sgo__n47050;
wire CLOCK_sgo__n47051;
wire CLOCK_slo__sro_n49350;
wire CLOCK_sgo__n47054;
wire CLOCK_slo__sro_n49382;
wire CLOCK_slo__sro_n49383;
wire CLOCK_slo__sro_n49384;
wire CLOCK_slo__sro_n51093;
wire CLOCK_slo__sro_n49386;
wire CLOCK_slo__sro_n49403;
wire CLOCK_opt_ipo_n46133;
wire CLOCK_slo__sro_n49426;
wire CLOCK_opt_ipo_n46137;
wire CLOCK_slo__sro_n49428;
wire CLOCK_slo__sro_n49429;
wire opt_ipo_n45556;
wire CLOCK_opt_ipo_n46146;
wire CLOCK_slo__sro_n49663;
wire CLOCK_slo__sro_n49664;
wire opt_ipo_n25394;
wire CLOCK_slo__sro_n49674;
wire CLOCK_slo__sro_n49713;
wire CLOCK_slo__sro_n49714;
wire CLOCK_slo__sro_n49726;
wire CLOCK_slo__sro_n61785;
wire CLOCK_slo__sro_n49727;
wire CLOCK_slo__sro_n49728;
wire CLOCK_slo__sro_n49758;
wire CLOCK_slo__sro_n61697;
wire CLOCK_slo__sro_n49759;
wire CLOCK_slo__sro_n49760;
wire CLOCK_slo__sro_n49761;
wire CLOCK_opt_ipo_n46189;
wire CLOCK_slo__sro_n49774;
wire CLOCK_slo__sro_n49775;
wire CLOCK_slo__sro_n49863;
wire CLOCK_slo__sro_n49864;
wire opt_ipo_n44394;
wire CLOCK_slo___n65042;
wire CLOCK_slo__sro_n49911;
wire CLOCK_slo__sro_n49912;
wire CLOCK_slo__sro_n49913;
wire CLOCK_slo__sro_n49937;
wire CLOCK_slo__sro_n49938;
wire CLOCK_slo__sro_n49939;
wire CLOCK_slo__sro_n49961;
wire CLOCK_slo__sro_n49962;
wire CLOCK_slo__sro_n50082;
wire CLOCK_slo__sro_n50068;
wire CLOCK_slo__sro_n50069;
wire CLOCK_slo__sro_n50070;
wire CLOCK_slo__sro_n50071;
wire CLOCK_slo__sro_n50097;
wire CLOCK_slo__sro_n50098;
wire CLOCK_slo__sro_n50131;
wire CLOCK_slo__sro_n50138;
wire CLOCK_slo__sro_n50139;
wire CLOCK_slo__sro_n50140;
wire CLOCK_slo__sro_n50141;
wire CLOCK_slo__sro_n50187;
wire CLOCK_slo__sro_n50188;
wire CLOCK_slo__sro_n50224;
wire CLOCK_slo__sro_n50225;
wire CLOCK_slo__sro_n50226;
wire CLOCK_opt_ipo_n46265;
wire CLOCK_slo__sro_n50227;
wire CLOCK_slo__sro_n50301;
wire CLOCK_slo__sro_n50302;
wire CLOCK_slo__sro_n50303;
wire CLOCK_slo__sro_n50319;
wire CLOCK_slo__sro_n50320;
wire CLOCK_slo__sro_n50321;
wire CLOCK_slo__sro_n50330;
wire CLOCK_slo__sro_n50331;
wire CLOCK_slo__sro_n50332;
wire CLOCK_slo__sro_n50362;
wire CLOCK_sgo__sro_n47110;
wire CLOCK_slo__sro_n50364;
wire CLOCK_slo__sro_n50400;
wire CLOCK_slo__sro_n50401;
wire CLOCK_slo__sro_n50402;
wire CLOCK_slo__sro_n50403;
wire CLOCK_slo__n50420;
wire CLOCK_slo__n50421;
wire CLOCK_slo__sro_n50433;
wire CLOCK_slo__sro_n65091;
wire CLOCK_slo__sro_n50547;
wire CLOCK_slo__sro_n50484;
wire CLOCK_slo__sro_n50522;
wire CLOCK_slo__sro_n50523;
wire CLOCK_slo__sro_n50524;
wire CLOCK_slo__sro_n50525;
wire CLOCK_slo__sro_n50657;
wire CLOCK_slo__sro_n50608;
wire CLOCK_slo__sro_n50609;
wire CLOCK_slo__sro_n50610;
wire CLOCK_slo__sro_n50611;
wire CLOCK_slo__sro_n50659;
wire CLOCK_slo__sro_n50660;
wire CLOCK_slo__sro_n50682;
wire CLOCK_slo__sro_n50730;
wire CLOCK_slo__sro_n50731;
wire CLOCK_slo__sro_n50793;
wire CLOCK_slo__sro_n50794;
wire CLOCK_slo__sro_n50830;
wire CLOCK_slo__sro_n50831;
wire CLOCK_slo__sro_n62824;
wire CLOCK_slo__sro_n50840;
wire CLOCK_slo__sro_n50841;
wire CLOCK_slo__sro_n50850;
wire CLOCK_slo__sro_n50862;
wire CLOCK_slo__sro_n50863;
wire CLOCK_slo__sro_n50864;
wire CLOCK_slo__sro_n50912;
wire CLOCK_slo__sro_n50913;
wire CLOCK_slo__n50956;
wire CLOCK_slo__sro_n50975;
wire CLOCK_slo__sro_n50976;
wire CLOCK_slo__sro_n50986;
wire CLOCK_slo__sro_n50987;
wire CLOCK_slo__sro_n51060;
wire CLOCK_slo__sro_n51061;
wire CLOCK_slo__sro_n51062;
wire opt_ipo_n44599;
wire CLOCK_slo__sro_n51094;
wire CLOCK_slo__sro_n51095;
wire CLOCK_slo__sro_n51133;
wire CLOCK_slo__sro_n51262;
wire CLOCK_slo__sro_n51306;
wire CLOCK_slo__sro_n51307;
wire CLOCK_slo__sro_n51308;
wire CLOCK_slo__sro_n51309;
wire CLOCK_slo__mro_n51372;
wire CLOCK_slo__mro_n51373;
wire CLOCK_slo__sro_n51475;
wire CLOCK_slo__sro_n51439;
wire CLOCK_slo__sro_n51440;
wire CLOCK_slo__sro_n51441;
wire CLOCK_slo__sro_n51442;
wire CLOCK_slo__mro_n51497;
wire CLOCK_slo__sro_n51513;
wire CLOCK_slo__mro_n51529;
wire CLOCK_slo__sro_n51542;
wire CLOCK_slo__sro_n51543;
wire CLOCK_slo__sro_n51544;
wire CLOCK_slo__sro_n51601;
wire CLOCK_slo__sro_n51602;
wire CLOCK_slo__sro_n51603;
wire CLOCK_slo__sro_n51604;
wire CLOCK_sgo__sro_n47109;
wire CLOCK_slo__sro_n51621;
wire CLOCK_slo__sro_n63269;
wire CLOCK_slo__sro_n51643;
wire CLOCK_slo__sro_n51644;
wire CLOCK_slo__sro_n51645;
wire CLOCK_slo__sro_n51724;
wire CLOCK_slo__sro_n53932;
wire CLOCK_slo__sro_n51725;
wire CLOCK_slo__sro_n51766;
wire CLOCK_slo__sro_n51773;
wire CLOCK_slo__sro_n51774;
wire CLOCK_slo__sro_n51775;
wire CLOCK_slo__sro_n51776;
wire CLOCK_slo__sro_n51853;
wire CLOCK_slo__sro_n51885;
wire CLOCK_slo__sro_n51886;
wire CLOCK_slo__sro_n51834;
wire CLOCK_slo__sro_n51835;
wire CLOCK_slo__sro_n51836;
wire CLOCK_slo__sro_n51887;
wire CLOCK_slo__sro_n51958;
wire CLOCK_slo__sro_n51959;
wire CLOCK_slo__sro_n51980;
wire CLOCK_slo__sro_n51981;
wire CLOCK_slo__sro_n51982;
wire CLOCK_slo__sro_n52124;
wire CLOCK_slo__sro_n52125;
wire CLOCK_slo__sro_n52126;
wire CLOCK_slo__sro_n52137;
wire CLOCK_slo__sro_n52054;
wire CLOCK_slo__sro_n52055;
wire CLOCK_slo__sro_n52056;
wire CLOCK_slo__sro_n52138;
wire CLOCK_slo__mro_n52164;
wire CLOCK_slo__mro_n52173;
wire CLOCK_slo__mro_n52174;
wire CLOCK_slo___n52225;
wire CLOCK_slo__sro_n52592;
wire CLOCK_slo__sro_n52593;
wire CLOCK_slo__sro_n52568;
wire CLOCK_slo__sro_n52569;
wire CLOCK_slo__sro_n52570;
wire CLOCK_slo__sro_n52540;
wire CLOCK_slo__sro_n52541;
wire CLOCK_slo__sro_n52542;
wire CLOCK_slo__sro_n52571;
wire CLOCK_slo__sro_n52595;
wire CLOCK_slo__sro_n52671;
wire CLOCK_slo__sro_n52915;
wire CLOCK_slo__sro_n52632;
wire CLOCK_slo__sro_n52633;
wire CLOCK_slo__sro_n52917;
wire CLOCK_slo__sro_n53419;
wire CLOCK_slo__sro_n52466;
wire CLOCK_slo__sro_n52635;
wire CLOCK_slo__sro_n52971;
wire CLOCK_slo__sro_n52972;
wire CLOCK_slo__sro_n53078;
wire CLOCK_slo__sro_n53079;
wire CLOCK_slo__sro_n53015;
wire CLOCK_slo__sro_n53339;
wire CLOCK_slo__sro_n52794;
wire CLOCK_slo__sro_n52795;
wire CLOCK_slo__sro_n53277;
wire CLOCK_slo__sro_n53278;
wire CLOCK_slo__sro_n53257;
wire CLOCK_slo__sro_n53064;
wire CLOCK_slo__sro_n53156;
wire CLOCK_slo__sro_n53157;
wire CLOCK_slo__sro_n53158;
wire CLOCK_slo__sro_n53159;
wire CLOCK_slo__sro_n53196;
wire CLOCK_slo__sro_n53197;
wire CLOCK_slo__sro_n53198;
wire CLOCK_slo__sro_n53406;
wire CLOCK_slo__sro_n53571;
wire CLOCK_slo__sro_n53258;
wire CLOCK_slo__sro_n53259;
wire CLOCK_slo__sro_n53260;
wire CLOCK_slo__n53562;
wire CLOCK_slo__sro_n53572;
wire CLOCK_slo__sro_n54099;
wire CLOCK_slo___n53904;
wire CLOCK_slo__n53697;
wire CLOCK_slo__sro_n54312;
wire CLOCK_slo__sro_n54100;
wire CLOCK_slo__sro_n54053;
wire CLOCK_slo__sro_n54054;
wire CLOCK_slo__sro_n53823;
wire CLOCK_slo__sro_n53824;
wire CLOCK_slo__sro_n53825;
wire CLOCK_slo__sro_n54055;
wire CLOCK_slo__sro_n53931;
wire CLOCK_slo__sro_n53892;
wire CLOCK_slo__sro_n53893;
wire CLOCK_slo__sro_n53894;
wire CLOCK_slo__n54187;
wire CLOCK_slo__n54289;
wire CLOCK_slo__sro_n54281;
wire CLOCK_slo__sro_n54313;
wire CLOCK_slo__sro_n54282;
wire CLOCK_slo__n54298;
wire CLOCK_slo__sro_n54314;
wire CLOCK_slo__sro_n54315;
wire CLOCK_slo__sro_n54488;
wire CLOCK_slo__sro_n54471;
wire CLOCK_slo__sro_n54472;
wire CLOCK_slo__sro_n54473;
wire CLOCK_slo__sro_n54474;
wire CLOCK_slo__sro_n54568;
wire CLOCK_slo__sro_n54569;
wire CLOCK_slo___n54911;
wire CLOCK_slo__sro_n54605;
wire CLOCK_slo__sro_n54698;
wire CLOCK_slo__sro_n54551;
wire CLOCK_slo__sro_n54552;
wire CLOCK_slo__sro_n54553;
wire CLOCK_slo__sro_n54554;
wire CLOCK_slo__n54674;
wire CLOCK_slo__sro_n54707;
wire CLOCK_slo__sro_n55060;
wire CLOCK_slo__sro_n54884;
wire CLOCK_slo__sro_n54885;
wire CLOCK_slo__sro_n54886;
wire CLOCK_slo___n64878;
wire CLOCK_slo__sro_n55019;
wire CLOCK_slo__sro_n54789;
wire CLOCK_slo__n55041;
wire CLOCK_slo__sro_n55020;
wire CLOCK_slo__sro_n54952;
wire CLOCK_slo__n54964;
wire CLOCK_slo__sro_n55021;
wire CLOCK_slo__sro_n55022;
wire CLOCK_slo__sro_n55023;
wire CLOCK_slo__sro_n55085;
wire CLOCK_slo__sro_n55086;
wire CLOCK_slo__sro_n55087;
wire CLOCK_slo__sro_n55103;
wire CLOCK_slo__sro_n55104;
wire CLOCK_slo__sro_n55105;
wire CLOCK_slo__sro_n55169;
wire CLOCK_slo__sro_n55156;
wire CLOCK_slo__sro_n55157;
wire CLOCK_slo__sro_n64272;
wire CLOCK_slo__sro_n55170;
wire CLOCK_slo__sro_n55171;
wire CLOCK_slo__n55377;
wire CLOCK_slo__sro_n55808;
wire CLOCK_slo__n55511;
wire CLOCK_slo__n55232;
wire CLOCK_slo__n55312;
wire CLOCK_slo__n55755;
wire CLOCK_slo__sro_n55400;
wire CLOCK_slo__sro_n55398;
wire CLOCK_slo__sro_n55399;
wire CLOCK_slo__n55465;
wire CLOCK_slo__n55647;
wire CLOCK_slo__n55658;
wire CLOCK_slo__sro_n55447;
wire CLOCK_slo__sro_n55448;
wire CLOCK_slo__sro_n55449;
wire CLOCK_slo__sro_n55810;
wire CLOCK_slo__n55860;
wire CLOCK_slo__n55865;
wire CLOCK_slo__sro_n55888;
wire CLOCK_slo__sro_n55889;
wire CLOCK_slo__sro_n55890;
wire CLOCK_slo__sro_n55784;
wire CLOCK_slo__sro_n55785;
wire CLOCK_slo__n55908;
wire CLOCK_slo__sro_n55930;
wire CLOCK_slo__sro_n56009;
wire CLOCK_slo__sro_n55959;
wire CLOCK_slo__sro_n56017;
wire CLOCK_slo__sro_n56018;
wire CLOCK_slo__sro_n56019;
wire CLOCK_slo__sro_n56057;
wire CLOCK_slo__sro_n56058;
wire CLOCK_slo__sro_n56059;
wire CLOCK_slo__sro_n56060;
wire CLOCK_slo__sro_n56037;
wire CLOCK_slo__n56237;
wire CLOCK_slo__n56232;
wire CLOCK_slo__sro_n56126;
wire CLOCK_slo__sro_n56306;
wire CLOCK_slo__sro_n56260;
wire CLOCK_slo__sro_n56261;
wire CLOCK_slo__sro_n56376;
wire CLOCK_slo__n56313;
wire CLOCK_slo__sro_n56377;
wire CLOCK_slo__sro_n56378;
wire CLOCK_slo__sro_n56379;
wire CLOCK_slo__n56418;
wire CLOCK_slo__sro_n56597;
wire CLOCK_slo__sro_n56598;
wire CLOCK_slo__sro_n56609;
wire CLOCK_slo__sro_n56610;
wire CLOCK_slo__n56713;
wire CLOCK_slo__n56467;
wire CLOCK_slo__sro_n56757;
wire CLOCK_slo__sro_n56895;
wire CLOCK_slo__sro_n56896;
wire CLOCK_slo__n57308;
wire CLOCK_slo__n56734;
wire CLOCK_slo__n56953;
wire CLOCK_slo__n56881;
wire CLOCK_slo__n56933;
wire CLOCK_slo__n56946;
wire CLOCK_slo__sro_n57154;
wire CLOCK_slo__sro_n57155;
wire CLOCK_slo__xsl_n57029;
wire CLOCK_slo__sro_n57132;
wire CLOCK_slo__n57242;
wire CLOCK_slo__sro_n57490;
wire CLOCK_slo__n57456;
wire CLOCK_slo__sro_n57699;
wire CLOCK_slo__n57518;
wire CLOCK_slo__n57483;
wire CLOCK_slo__n57523;
wire CLOCK_slo__sro_n57700;
wire CLOCK_slo__n57534;
wire CLOCK_slo__n57556;
wire CLOCK_slo___n57806;
wire CLOCK_slo__n57547;
wire CLOCK_slo__sro_n57701;
wire CLOCK_slo__sro_n57685;
wire CLOCK_slo__sro_n57686;
wire CLOCK_slo__sro_n57687;
wire CLOCK_slo__n57906;
wire CLOCK_slo__n57799;
wire CLOCK_slo__n57760;
wire CLOCK_slo__n57977;
wire CLOCK_slo__n57899;
wire CLOCK_slo__n57874;
wire CLOCK_slo__sro_n58451;
wire CLOCK_slo__n57743;
wire CLOCK_slo__n58182;
wire CLOCK_slo__n58099;
wire CLOCK_slo__sro_n58144;
wire CLOCK_slo__sro_n58145;
wire CLOCK_slo__sro_n58146;
wire CLOCK_slo__sro_n58465;
wire CLOCK_slo__n58195;
wire CLOCK_slo__sro_n58342;
wire CLOCK_slo__sro_n58313;
wire CLOCK_slo__sro_n58314;
wire CLOCK_slo__sro_n58234;
wire CLOCK_slo__sro_n58235;
wire CLOCK_slo__sro_n58315;
wire CLOCK_slo__sro_n58708;
wire CLOCK_slo__n58422;
wire CLOCK_slo___n58400;
wire CLOCK_slo__sro_n58709;
wire CLOCK_slo__sro_n58698;
wire spw__n66802;
wire CLOCK_slo__sro_n58611;
wire CLOCK_slo__sro_n58699;
wire CLOCK_slo__sro_n58700;
wire CLOCK_slo__sro_n58710;
wire CLOCK_slo__sro_n58765;
wire CLOCK_slo__sro_n58518;
wire CLOCK_slo__sro_n58519;
wire CLOCK_slo__sro_n58520;
wire CLOCK_slo__sro_n58521;
wire CLOCK_slo__sro_n58766;
wire CLOCK_slo__sro_n58846;
wire CLOCK_slo__sro_n58847;
wire CLOCK_slo__sro_n58904;
wire CLOCK_slo__sro_n58905;
wire CLOCK_slo__sro_n58906;
wire CLOCK_slo__sro_n58907;
wire CLOCK_slo__sro_n59280;
wire CLOCK_slo__sro_n59281;
wire CLOCK_slo__sro_n59126;
wire CLOCK_slo__sro_n59056;
wire CLOCK_slo__sro_n59057;
wire CLOCK_slo__sro_n59058;
wire CLOCK_slo__sro_n59127;
wire CLOCK_slo__sro_n59128;
wire CLOCK_slo__sro_n62893;
wire CLOCK_slo__sro_n59283;
wire CLOCK_slo__sro_n59303;
wire CLOCK_slo__sro_n59027;
wire CLOCK_slo__sro_n59028;
wire CLOCK_slo__sro_n59029;
wire CLOCK_slo__sro_n63004;
wire CLOCK_slo__sro_n59343;
wire CLOCK_slo__sro_n59344;
wire CLOCK_slo__sro_n59345;
wire CLOCK_slo__sro_n59447;
wire CLOCK_slo__sro_n59448;
wire CLOCK_slo__sro_n59468;
wire CLOCK_slo__sro_n59469;
wire CLOCK_slo__sro_n59533;
wire CLOCK_slo__sro_n59534;
wire CLOCK_slo__sro_n59535;
wire CLOCK_slo__sro_n59549;
wire CLOCK_slo__sro_n59550;
wire CLOCK_slo__sro_n59551;
wire CLOCK_slo__sro_n59728;
wire CLOCK_slo__sro_n59712;
wire CLOCK_slo__sro_n59713;
wire CLOCK_slo__sro_n59714;
wire CLOCK_slo__sro_n59730;
wire CLOCK_slo__sro_n59951;
wire CLOCK_slo__sro_n59961;
wire CLOCK_slo__sro_n59962;
wire CLOCK_slo__sro_n60053;
wire CLOCK_slo__sro_n60054;
wire CLOCK_slo__sro_n59842;
wire CLOCK_slo__sro_n59843;
wire CLOCK_slo__sro_n59773;
wire CLOCK_slo__sro_n59774;
wire CLOCK_slo__sro_n59775;
wire CLOCK_slo__sro_n59845;
wire CLOCK_slo__sro_n60126;
wire CLOCK_slo__sro_n60127;
wire CLOCK_slo__sro_n60276;
wire CLOCK_slo__sro_n60277;
wire CLOCK_slo__sro_n60278;
wire CLOCK_slo__sro_n60309;
wire CLOCK_slo__sro_n60310;
wire CLOCK_slo__n60587;
wire CLOCK_slo__sro_n60604;
wire CLOCK_slo__sro_n60605;
wire CLOCK_slo__sro_n60639;
wire CLOCK_slo__sro_n60640;
wire CLOCK_slo__sro_n60641;
wire CLOCK_slo__sro_n60642;
wire CLOCK_slo__sro_n60680;
wire CLOCK_slo__sro_n60681;
wire CLOCK_slo__sro_n60763;
wire CLOCK_slo__sro_n60777;
wire CLOCK_slo__sro_n60778;
wire CLOCK_slo__sro_n60812;
wire CLOCK_slo__sro_n60813;
wire CLOCK_slo__sro_n60814;
wire CLOCK_slo__sro_n60815;


INV_X1 i_0_0_154 (.ZN (n_0_0_28), .A (Multiplier[31]));
BUF_X1 CLOCK_sgo__L2_c2_c51290 (.Z (n_6_1_874), .A (CLOCK_sgo__n47093));
INV_X2 i_0_0_152 (.ZN (n_0_0_26), .A (n_0_61));
NOR4_X1 i_0_0_151 (.ZN (n_0_0_25), .A1 (Multiplicand[15]), .A2 (Multiplicand[10])
    , .A3 (Multiplicand[9]), .A4 (Multiplicand[8]));
NOR4_X1 i_0_0_150 (.ZN (n_0_0_24), .A1 (Multiplicand[14]), .A2 (Multiplicand[13])
    , .A3 (Multiplicand[12]), .A4 (Multiplicand[11]));
NOR4_X1 i_0_0_149 (.ZN (n_0_0_23), .A1 (Multiplicand[7]), .A2 (Multiplicand[2]), .A3 (Multiplicand[1]), .A4 (Multiplicand[0]));
NOR4_X1 i_0_0_148 (.ZN (n_0_0_22), .A1 (Multiplicand[6]), .A2 (Multiplicand[5]), .A3 (Multiplicand[4]), .A4 (Multiplicand[3]));
NAND4_X1 i_0_0_147 (.ZN (n_0_0_21), .A1 (n_0_0_25), .A2 (n_0_0_24), .A3 (n_0_0_23), .A4 (n_0_0_22));
NOR4_X1 i_0_0_146 (.ZN (n_0_0_20), .A1 (Multiplicand[27]), .A2 (Multiplicand[26])
    , .A3 (Multiplicand[25]), .A4 (Multiplicand[16]));
NOR4_X1 i_0_0_145 (.ZN (n_0_0_19), .A1 (Multiplicand[31]), .A2 (Multiplicand[30])
    , .A3 (Multiplicand[29]), .A4 (Multiplicand[28]));
NOR4_X1 i_0_0_144 (.ZN (n_0_0_18), .A1 (Multiplicand[24]), .A2 (Multiplicand[19])
    , .A3 (Multiplicand[18]), .A4 (Multiplicand[17]));
NOR4_X1 i_0_0_143 (.ZN (n_0_0_17), .A1 (Multiplicand[23]), .A2 (Multiplicand[22])
    , .A3 (Multiplicand[21]), .A4 (Multiplicand[20]));
NAND4_X1 i_0_0_142 (.ZN (n_0_0_16), .A1 (n_0_0_20), .A2 (n_0_0_19), .A3 (n_0_0_18), .A4 (n_0_0_17));
NOR2_X1 i_0_0_141 (.ZN (n_0_0_15), .A1 (n_0_0_21), .A2 (n_0_0_16));
NOR4_X1 i_0_0_140 (.ZN (n_0_0_14), .A1 (drc_ipoPP_7), .A2 (drc_ipoPP_6), .A3 (Multiplier[25]), .A4 (Multiplier[24]));
NOR4_X1 i_0_0_139 (.ZN (n_0_0_13), .A1 (hfn_ipo_n26), .A2 (drc_ipo_n26625), .A3 (drc_ipo_n26624), .A4 (sgo__n1276));
NOR4_X1 i_0_0_138 (.ZN (n_0_0_12), .A1 (drc_ipoPP_5), .A2 (drc_ipo_n26614), .A3 (drc_ipo_n26613), .A4 (drc_ipoPP_4));
NOR4_X1 i_0_0_137 (.ZN (n_0_0_11), .A1 (Multiplier[22]), .A2 (drc_ipo_n26616), .A3 (Multiplier[20]), .A4 (drc_ipoPP_3));
NAND4_X1 i_0_0_136 (.ZN (n_0_0_10), .A1 (n_0_0_14), .A2 (n_0_0_13), .A3 (n_0_0_12), .A4 (n_0_0_11));
NOR4_X1 i_0_0_135 (.ZN (n_0_0_9), .A1 (Multiplier[7]), .A2 (slo__n3804), .A3 (sgo__n1306), .A4 (slo__n18930));
NOR4_X1 i_0_0_134 (.ZN (n_0_0_8), .A1 (drc_ipo_n26610), .A2 (slo__n11938), .A3 (slo__n4958), .A4 (slo__n4944));
NOR4_X1 i_0_0_133 (.ZN (n_0_0_7), .A1 (Multiplier[11]), .A2 (Multiplier[10]), .A3 (Multiplier[9]), .A4 (Multiplier[8]));
NOR3_X1 i_0_0_132 (.ZN (n_0_0_6), .A1 (Multiplier[14]), .A2 (Multiplier[13]), .A3 (Multiplier[12]));
NAND4_X1 i_0_0_131 (.ZN (n_0_0_5), .A1 (n_0_0_9), .A2 (n_0_0_8), .A3 (n_0_0_7), .A4 (n_0_0_6));
OR2_X1 i_0_0_130 (.ZN (n_0_0_4), .A1 (n_0_0_10), .A2 (n_0_0_5));
INV_X1 i_0_0_129 (.ZN (n_0_0_3), .A (n_0_0_4));
AOI21_X1 i_0_0_128 (.ZN (n_0_0_2), .A (n_0_0_15), .B1 (n_0_0_3), .B2 (n_0_0_28));
AND2_X4 i_0_0_127 (.ZN (n_0_124), .A1 (opt_ipo_n23872), .A2 (hfn_ipo_n35));
NAND2_X1 CLOCK_slo__sro_c68586 (.ZN (CLOCK_slo__sro_n61786), .A1 (n_6_2051), .A2 (n_6_1_133));
AOI21_X4 slo__sro_c16778 (.ZN (slo__sro_n15079), .A (sgo__sro_n1676), .B1 (n_6_35), .B2 (n_6_1_1114));
AND2_X4 i_0_0_123 (.ZN (n_0_120), .A1 (CLOCK_opt_ipo_n45736), .A2 (hfn_ipo_n35));
AND2_X2 i_0_0_122 (.ZN (n_0_119), .A1 (n_57), .A2 (hfn_ipo_n35));
AND2_X2 i_0_0_121 (.ZN (n_0_118), .A1 (n_56), .A2 (hfn_ipo_n35));
AND2_X1 i_0_0_120 (.ZN (n_0_117), .A1 (n_55), .A2 (hfn_ipo_n35));
AND2_X1 i_0_0_119 (.ZN (n_0_116), .A1 (n_54), .A2 (hfn_ipo_n35));
AND2_X2 i_0_0_118 (.ZN (n_0_115), .A1 (n_6_1_52), .A2 (hfn_ipo_n35));
AND2_X1 i_0_0_117 (.ZN (n_0_114), .A1 (n_52), .A2 (hfn_ipo_n35));
AND2_X1 i_0_0_116 (.ZN (n_0_113), .A1 (n_51), .A2 (hfn_ipo_n35));
AND2_X1 i_0_0_115 (.ZN (n_0_112), .A1 (n_50), .A2 (hfn_ipo_n35));
AND2_X2 i_0_0_114 (.ZN (n_0_111), .A1 (n_49), .A2 (hfn_ipo_n35));
AND2_X4 i_0_0_113 (.ZN (n_0_110), .A1 (n_48), .A2 (hfn_ipo_n35));
AND2_X1 i_0_0_112 (.ZN (n_0_109), .A1 (n_47), .A2 (hfn_ipo_n35));
AND2_X1 i_0_0_111 (.ZN (n_0_108), .A1 (n_46), .A2 (hfn_ipo_n35));
AND2_X2 i_0_0_110 (.ZN (n_0_107), .A1 (n_45), .A2 (hfn_ipo_n35));
AND2_X1 i_0_0_109 (.ZN (n_0_106), .A1 (n_44), .A2 (hfn_ipo_n35));
AND2_X1 i_0_0_108 (.ZN (n_0_105), .A1 (n_43), .A2 (hfn_ipo_n35));
AND2_X1 i_0_0_107 (.ZN (n_0_104), .A1 (n_42), .A2 (hfn_ipo_n35));
AND2_X4 i_0_0_106 (.ZN (n_0_103), .A1 (n_41), .A2 (hfn_ipo_n35));
AND2_X1 i_0_0_105 (.ZN (n_0_102), .A1 (n_40), .A2 (hfn_ipo_n35));
AND2_X2 i_0_0_104 (.ZN (n_0_101), .A1 (n_39), .A2 (hfn_ipo_n35));
AND2_X1 i_0_0_103 (.ZN (n_0_100), .A1 (n_38), .A2 (hfn_ipo_n35));
AND2_X2 i_0_0_102 (.ZN (n_0_99), .A1 (n_37), .A2 (hfn_ipo_n35));
AND2_X1 i_0_0_101 (.ZN (n_0_98), .A1 (n_36), .A2 (hfn_ipo_n35));
AND2_X1 i_0_0_100 (.ZN (n_0_97), .A1 (n_35), .A2 (hfn_ipo_n35));
AND2_X2 i_0_0_99 (.ZN (n_0_96), .A1 (n_34), .A2 (hfn_ipo_n35));
AND2_X1 i_0_0_98 (.ZN (n_0_95), .A1 (n_33), .A2 (hfn_ipo_n35));
AND2_X1 i_0_0_97 (.ZN (n_0_94), .A1 (n_32), .A2 (hfn_ipo_n35));
AND2_X1 i_0_0_96 (.ZN (n_0_93), .A1 (n_31), .A2 (hfn_ipo_n35));
AND2_X1 i_0_0_95 (.ZN (n_0_92), .A1 (n_30), .A2 (hfn_ipo_n35));
AND2_X1 i_0_0_94 (.ZN (n_0_91), .A1 (n_29), .A2 (hfn_ipo_n36));
AND2_X2 i_0_0_93 (.ZN (n_0_90), .A1 (n_28), .A2 (hfn_ipo_n36));
AND2_X1 i_0_0_92 (.ZN (n_0_89), .A1 (n_27), .A2 (hfn_ipo_n36));
AND2_X2 i_0_0_91 (.ZN (n_0_88), .A1 (n_26), .A2 (hfn_ipo_n36));
AND2_X1 i_0_0_90 (.ZN (n_0_87), .A1 (n_25), .A2 (hfn_ipo_n36));
AND2_X1 i_0_0_89 (.ZN (n_0_86), .A1 (n_24), .A2 (hfn_ipo_n36));
AND2_X1 i_0_0_88 (.ZN (n_0_85), .A1 (n_23), .A2 (hfn_ipo_n36));
AND2_X2 i_0_0_87 (.ZN (n_0_84), .A1 (n_22), .A2 (hfn_ipo_n36));
AND2_X1 i_0_0_86 (.ZN (n_0_83), .A1 (n_21), .A2 (hfn_ipo_n36));
AND2_X1 i_0_0_85 (.ZN (n_0_82), .A1 (n_20), .A2 (hfn_ipo_n36));
AND2_X1 i_0_0_84 (.ZN (n_0_81), .A1 (n_19), .A2 (hfn_ipo_n36));
AND2_X1 i_0_0_83 (.ZN (n_0_80), .A1 (n_18), .A2 (hfn_ipo_n36));
AND2_X1 i_0_0_82 (.ZN (n_0_79), .A1 (n_17), .A2 (hfn_ipo_n36));
AND2_X1 i_0_0_81 (.ZN (n_0_78), .A1 (n_16), .A2 (hfn_ipo_n36));
AND2_X2 i_0_0_80 (.ZN (n_0_77), .A1 (n_15), .A2 (hfn_ipo_n36));
AND2_X1 i_0_0_79 (.ZN (n_0_76), .A1 (n_14), .A2 (hfn_ipo_n36));
AND2_X1 i_0_0_78 (.ZN (n_0_75), .A1 (n_13), .A2 (hfn_ipo_n36));
AND2_X1 i_0_0_77 (.ZN (n_0_74), .A1 (n_12), .A2 (hfn_ipo_n36));
AND2_X1 i_0_0_76 (.ZN (n_0_73), .A1 (n_11), .A2 (hfn_ipo_n36));
AND2_X1 i_0_0_75 (.ZN (n_0_72), .A1 (n_10), .A2 (hfn_ipo_n36));
AND2_X1 i_0_0_74 (.ZN (n_0_71), .A1 (n_9), .A2 (hfn_ipo_n36));
AND2_X1 i_0_0_73 (.ZN (n_0_70), .A1 (n_8), .A2 (hfn_ipo_n36));
AND2_X1 i_0_0_72 (.ZN (n_0_69), .A1 (n_7), .A2 (hfn_ipo_n36));
AND2_X1 i_0_0_71 (.ZN (n_0_68), .A1 (n_6), .A2 (hfn_ipo_n36));
AND2_X1 i_0_0_70 (.ZN (n_0_67), .A1 (n_5), .A2 (hfn_ipo_n36));
AND2_X1 i_0_0_69 (.ZN (n_0_66), .A1 (n_4), .A2 (hfn_ipo_n36));
AND2_X1 i_0_0_68 (.ZN (n_0_65), .A1 (n_3), .A2 (hfn_ipo_n36));
AND2_X1 i_0_0_67 (.ZN (n_0_64), .A1 (n_2), .A2 (hfn_ipo_n36));
AND2_X1 i_0_0_66 (.ZN (n_0_63), .A1 (n_1), .A2 (hfn_ipo_n36));
AND2_X1 i_0_0_65 (.ZN (Product[0]), .A1 (n_0), .A2 (hfn_ipo_n36));
NAND2_X1 i_0_0_64 (.ZN (n_0_0_1), .A1 (Multiplier[31]), .A2 (n_0_0_3));
NAND2_X1 i_0_0_63 (.ZN (n_0_0_0), .A1 (n_0_124), .A2 (hfn_ipo_n33));
OAI21_X2 i_0_0_62 (.ZN (Product[63]), .A (n_0_0_0), .B1 (opt_ipo_n43864), .B2 (hfn_ipo_n33));
OAI21_X4 i_0_0_61 (.ZN (Product[62]), .A (n_0_0_0), .B1 (n_0_0_26), .B2 (hfn_ipo_n33));
MUX2_X1 i_0_0_60 (.Z (Product[61]), .A (n_0_60), .B (slo__mro_n33266), .S (hfn_ipo_n33));
AOI21_X1 slo__sro_c44166 (.ZN (slo__sro_n6737), .A (slo__sro_n39795), .B1 (n_6_1837), .B2 (n_6_1_135));
MUX2_X1 i_0_0_58 (.Z (Product[59]), .A (n_0_58), .B (slo__sro_n14967), .S (hfn_ipo_n33));
MUX2_X1 i_0_0_57 (.Z (Product[58]), .A (n_0_57), .B (n_0_120), .S (hfn_ipo_n33));
MUX2_X1 i_0_0_56 (.Z (Product[57]), .A (n_0_56), .B (n_0_119), .S (hfn_ipo_n33));
MUX2_X1 i_0_0_55 (.Z (Product[56]), .A (n_0_55), .B (n_0_118), .S (hfn_ipo_n33));
MUX2_X1 i_0_0_54 (.Z (Product[55]), .A (n_0_54), .B (n_0_117), .S (hfn_ipo_n33));
MUX2_X1 i_0_0_53 (.Z (Product[54]), .A (n_0_53), .B (n_0_116), .S (hfn_ipo_n33));
MUX2_X1 i_0_0_52 (.Z (Product[53]), .A (n_0_52), .B (n_0_115), .S (hfn_ipo_n33));
MUX2_X1 i_0_0_51 (.Z (Product[52]), .A (n_0_51), .B (n_0_114), .S (hfn_ipo_n33));
MUX2_X1 i_0_0_50 (.Z (Product[51]), .A (n_0_50), .B (n_0_113), .S (hfn_ipo_n33));
MUX2_X1 i_0_0_49 (.Z (Product[50]), .A (n_0_49), .B (n_0_112), .S (hfn_ipo_n33));
MUX2_X1 i_0_0_48 (.Z (Product[49]), .A (n_0_48), .B (n_0_111), .S (hfn_ipo_n33));
MUX2_X1 i_0_0_47 (.Z (Product[48]), .A (n_0_47), .B (n_0_110), .S (hfn_ipo_n33));
MUX2_X1 i_0_0_46 (.Z (Product[47]), .A (n_0_46), .B (n_0_109), .S (hfn_ipo_n33));
MUX2_X1 i_0_0_45 (.Z (Product[46]), .A (n_0_45), .B (n_0_108), .S (hfn_ipo_n33));
MUX2_X1 i_0_0_44 (.Z (Product[45]), .A (n_0_44), .B (n_0_107), .S (hfn_ipo_n33));
MUX2_X1 i_0_0_43 (.Z (Product[44]), .A (n_0_43), .B (n_0_106), .S (hfn_ipo_n33));
MUX2_X1 i_0_0_42 (.Z (Product[43]), .A (n_0_42), .B (n_0_105), .S (hfn_ipo_n33));
MUX2_X1 i_0_0_41 (.Z (Product[42]), .A (n_0_41), .B (n_0_104), .S (hfn_ipo_n33));
MUX2_X1 i_0_0_40 (.Z (Product[41]), .A (n_0_40), .B (n_0_103), .S (hfn_ipo_n33));
MUX2_X1 i_0_0_39 (.Z (Product[40]), .A (n_0_39), .B (n_0_102), .S (hfn_ipo_n33));
MUX2_X1 i_0_0_38 (.Z (Product[39]), .A (n_0_38), .B (n_0_101), .S (hfn_ipo_n33));
MUX2_X1 i_0_0_37 (.Z (Product[38]), .A (n_0_37), .B (n_0_100), .S (hfn_ipo_n33));
MUX2_X2 i_0_0_36 (.Z (Product[37]), .A (n_0_36), .B (n_0_99), .S (hfn_ipo_n33));
MUX2_X1 i_0_0_35 (.Z (Product[36]), .A (n_0_35), .B (n_0_98), .S (hfn_ipo_n33));
MUX2_X1 i_0_0_34 (.Z (Product[35]), .A (n_0_34), .B (n_0_97), .S (hfn_ipo_n33));
MUX2_X1 i_0_0_33 (.Z (Product[34]), .A (n_0_33), .B (n_0_96), .S (hfn_ipo_n33));
MUX2_X1 i_0_0_32 (.Z (Product[33]), .A (n_0_32), .B (n_0_95), .S (hfn_ipo_n33));
MUX2_X1 i_0_0_31 (.Z (Product[32]), .A (n_0_31), .B (n_0_94), .S (hfn_ipo_n33));
MUX2_X1 i_0_0_30 (.Z (Product[31]), .A (n_0_30), .B (n_0_93), .S (hfn_ipo_n33));
MUX2_X1 i_0_0_29 (.Z (Product[30]), .A (n_0_29), .B (n_0_92), .S (hfn_ipo_n33));
MUX2_X1 i_0_0_28 (.Z (Product[29]), .A (n_0_28), .B (n_0_91), .S (hfn_ipo_n34));
MUX2_X1 i_0_0_27 (.Z (Product[28]), .A (n_0_27), .B (n_0_90), .S (hfn_ipo_n34));
MUX2_X1 i_0_0_26 (.Z (Product[27]), .A (n_0_26), .B (n_0_89), .S (hfn_ipo_n34));
MUX2_X1 i_0_0_25 (.Z (Product[26]), .A (n_0_25), .B (n_0_88), .S (hfn_ipo_n34));
MUX2_X1 i_0_0_24 (.Z (Product[25]), .A (n_0_24), .B (n_0_87), .S (hfn_ipo_n34));
MUX2_X1 i_0_0_23 (.Z (Product[24]), .A (n_0_23), .B (n_0_86), .S (hfn_ipo_n34));
MUX2_X1 i_0_0_22 (.Z (Product[23]), .A (n_0_22), .B (n_0_85), .S (hfn_ipo_n34));
MUX2_X1 i_0_0_21 (.Z (Product[22]), .A (n_0_21), .B (n_0_84), .S (hfn_ipo_n34));
MUX2_X1 i_0_0_20 (.Z (Product[21]), .A (n_0_20), .B (n_0_83), .S (hfn_ipo_n34));
MUX2_X1 i_0_0_19 (.Z (Product[20]), .A (n_0_19), .B (n_0_82), .S (hfn_ipo_n34));
MUX2_X1 i_0_0_18 (.Z (Product[19]), .A (n_0_18), .B (n_0_81), .S (hfn_ipo_n34));
MUX2_X1 i_0_0_17 (.Z (Product[18]), .A (n_0_17), .B (n_0_80), .S (hfn_ipo_n34));
MUX2_X1 i_0_0_16 (.Z (Product[17]), .A (n_0_16), .B (n_0_79), .S (hfn_ipo_n34));
MUX2_X1 i_0_0_15 (.Z (Product[16]), .A (n_0_15), .B (n_0_78), .S (hfn_ipo_n34));
MUX2_X1 i_0_0_14 (.Z (Product[15]), .A (n_0_14), .B (n_0_77), .S (hfn_ipo_n34));
MUX2_X2 i_0_0_13 (.Z (Product[14]), .A (n_0_13), .B (n_0_76), .S (hfn_ipo_n34));
MUX2_X1 i_0_0_12 (.Z (Product[13]), .A (n_0_12), .B (n_0_75), .S (hfn_ipo_n34));
MUX2_X1 i_0_0_11 (.Z (Product[12]), .A (n_0_11), .B (n_0_74), .S (hfn_ipo_n34));
MUX2_X1 i_0_0_10 (.Z (Product[11]), .A (n_0_10), .B (n_0_73), .S (hfn_ipo_n34));
MUX2_X1 i_0_0_9 (.Z (Product[10]), .A (n_0_9), .B (n_0_72), .S (hfn_ipo_n34));
MUX2_X1 i_0_0_8 (.Z (Product[9]), .A (n_0_8), .B (n_0_71), .S (hfn_ipo_n34));
MUX2_X1 i_0_0_7 (.Z (Product[8]), .A (n_0_7), .B (n_0_70), .S (hfn_ipo_n34));
MUX2_X1 i_0_0_6 (.Z (Product[7]), .A (n_0_6), .B (n_0_69), .S (hfn_ipo_n34));
MUX2_X1 i_0_0_5 (.Z (Product[6]), .A (n_0_5), .B (n_0_68), .S (hfn_ipo_n34));
MUX2_X1 i_0_0_4 (.Z (Product[5]), .A (n_0_4), .B (n_0_67), .S (hfn_ipo_n34));
MUX2_X1 i_0_0_3 (.Z (Product[4]), .A (n_0_3), .B (n_0_66), .S (hfn_ipo_n34));
MUX2_X1 i_0_0_2 (.Z (Product[3]), .A (n_0_2), .B (n_0_65), .S (hfn_ipo_n34));
MUX2_X1 i_0_0_1 (.Z (Product[2]), .A (n_0_1), .B (n_0_64), .S (hfn_ipo_n34));
MUX2_X1 i_0_0_0 (.Z (Product[1]), .A (n_0_0), .B (n_0_63), .S (hfn_ipo_n34));
datapath__0_253 i_0_4 (.p_1 ({n_0_62, n_0_61, n_0_60, n_0_59, n_0_58, n_0_57, n_0_56, 
    n_0_55, n_0_54, n_0_53, n_0_52, n_0_51, n_0_50, n_0_49, n_0_48, n_0_47, n_0_46, 
    n_0_45, n_0_44, n_0_43, n_0_42, n_0_41, n_0_40, n_0_39, n_0_38, n_0_37, n_0_36, 
    n_0_35, n_0_34, n_0_33, n_0_32, n_0_31, n_0_30, n_0_29, n_0_28, n_0_27, n_0_26, 
    n_0_25, n_0_24, n_0_23, n_0_22, n_0_21, n_0_20, n_0_19, n_0_18, n_0_17, n_0_16, 
    n_0_15, n_0_14, n_0_13, n_0_12, n_0_11, n_0_10, n_0_9, n_0_8, n_0_7, n_0_6, n_0_5, 
    n_0_4, n_0_3, n_0_2, n_0_1, n_0_0, uc_62}), .p_0 ({uc_61, n_0_124, slo__mro_n33266, 
    slo__mro_n33299, slo__sro_n14967, n_0_120, n_0_119, n_0_118, n_0_117, n_0_116, 
    n_0_115, n_0_114, n_0_113, n_0_112, n_0_111, n_0_110, n_0_109, n_0_108, n_0_107, 
    n_0_106, n_0_105, n_0_104, n_0_103, n_0_102, n_0_101, n_0_100, n_0_99, n_0_98, 
    n_0_97, n_0_96, n_0_95, n_0_94, n_0_93, n_0_92, n_0_91, n_0_90, n_0_89, n_0_88, 
    n_0_87, n_0_86, n_0_85, n_0_84, n_0_83, n_0_82, n_0_81, n_0_80, n_0_79, n_0_78, 
    n_0_77, n_0_76, n_0_75, n_0_74, n_0_73, n_0_72, n_0_71, n_0_70, n_0_69, n_0_68, 
    n_0_67, n_0_66, n_0_65, n_0_64, n_0_63, Product[0]}));
INV_X4 i_6_1_2139 (.ZN (n_6_1_1145), .A (Multiplicand[30]));
INV_X1 i_6_1_2138 (.ZN (n_6_1_1144), .A (Multiplicand[29]));
INV_X1 i_6_1_2137 (.ZN (n_6_1_1143), .A (Multiplicand[28]));
INV_X1 i_6_1_2136 (.ZN (n_6_1_1142), .A (Multiplicand[27]));
INV_X1 i_6_1_2135 (.ZN (n_6_1_1141), .A (Multiplicand[26]));
INV_X1 i_6_1_2134 (.ZN (n_6_1_1140), .A (Multiplicand[25]));
INV_X1 i_6_1_2133 (.ZN (n_6_1_1139), .A (Multiplicand[24]));
INV_X1 i_6_1_2132 (.ZN (n_6_1_1138), .A (Multiplicand[23]));
INV_X1 i_6_1_2131 (.ZN (n_6_1_1137), .A (Multiplicand[22]));
INV_X1 i_6_1_2130 (.ZN (n_6_1_1136), .A (Multiplicand[21]));
INV_X1 i_6_1_2129 (.ZN (n_6_1_1135), .A (Multiplicand[20]));
INV_X1 i_6_1_2128 (.ZN (n_6_1_1134), .A (Multiplicand[19]));
INV_X1 i_6_1_2127 (.ZN (n_6_1_1133), .A (Multiplicand[18]));
INV_X1 i_6_1_2126 (.ZN (n_6_1_1132), .A (Multiplicand[17]));
INV_X1 i_6_1_2125 (.ZN (n_6_1_1131), .A (Multiplicand[16]));
INV_X1 i_6_1_2124 (.ZN (n_6_1_1130), .A (Multiplicand[15]));
INV_X1 i_6_1_2123 (.ZN (n_6_1_1129), .A (Multiplicand[14]));
INV_X1 i_6_1_2122 (.ZN (n_6_1_1128), .A (Multiplicand[13]));
INV_X1 i_6_1_2121 (.ZN (n_6_1_1127), .A (Multiplicand[12]));
INV_X1 i_6_1_2120 (.ZN (n_6_1_1126), .A (Multiplicand[11]));
INV_X1 i_6_1_2119 (.ZN (n_6_1_1125), .A (Multiplicand[10]));
INV_X1 i_6_1_2118 (.ZN (n_6_1_1124), .A (Multiplicand[9]));
INV_X1 i_6_1_2117 (.ZN (n_6_1_1123), .A (Multiplicand[8]));
INV_X1 i_6_1_2116 (.ZN (n_6_1_1122), .A (Multiplicand[7]));
INV_X1 i_6_1_2115 (.ZN (n_6_1_1121), .A (Multiplicand[6]));
INV_X1 i_6_1_2114 (.ZN (n_6_1_1120), .A (Multiplicand[5]));
INV_X1 i_6_1_2113 (.ZN (n_6_1_1119), .A (Multiplicand[4]));
INV_X1 i_6_1_2112 (.ZN (n_6_1_1118), .A (Multiplicand[3]));
INV_X1 i_6_1_2111 (.ZN (n_6_1_1117), .A (Multiplicand[2]));
INV_X1 i_6_1_2110 (.ZN (n_6_1_1116), .A (Multiplicand[1]));
INV_X1 i_6_1_2109 (.ZN (n_6_1_1115), .A (Multiplicand[0]));
AND2_X1 i_6_1_2108 (.ZN (n_6_2913), .A1 (Multiplicand[0]), .A2 (n_6_30));
NOR2_X1 i_6_1_2107 (.ZN (sgo__n714), .A1 (Multiplicand[1]), .A2 (n_6_1_1115));
AOI22_X1 i_6_1_2106 (.ZN (n_6_1_1113), .A1 (n_6_62), .A2 (n_6_1_1114), .B1 (Multiplicand[1]), .B2 (n_6_30));
INV_X1 i_6_1_2105 (.ZN (n_6_2912), .A (n_6_1_1113));
NOR2_X2 i_6_1_2104 (.ZN (sgo__n711), .A1 (n_6_1_1116), .A2 (Multiplicand[0]));
NAND2_X1 slo__sro_c33833 (.ZN (slo__sro_n30286), .A1 (n_6_1099), .A2 (slo___n23277));
INV_X1 i_6_1_2102 (.ZN (n_6_2911), .A (n_6_1_1111));
NOR2_X2 i_6_1_2101 (.ZN (sgo__n691), .A1 (n_6_1_1116), .A2 (n_6_1_1115));
AOI222_X1 i_6_1_2100 (.ZN (n_6_1_1109), .A1 (hfn_ipo_n30), .A2 (opt_ipo_n24358), .B1 (n_6_28)
    , .B2 (slo__n30589), .C1 (n_6_60), .C2 (n_6_1_1114));
INV_X1 i_6_1_2099 (.ZN (n_6_2910), .A (n_6_1_1109));
BUF_X32 drc_ipo_c29958 (.Z (drc_ipo_n26581), .A (n_6_19));
INV_X1 i_6_1_2097 (.ZN (n_6_2909), .A (slo__sro_n2408));
AOI22_X1 slo__sro_c2348 (.ZN (slo__sro_n2401), .A1 (n_6_25), .A2 (opt_ipo_n24358)
    , .B1 (CLOCK_sgo__n47054), .B2 (slo__n30589));
INV_X1 i_6_1_2095 (.ZN (n_6_2908), .A (slo__sro_n2370));
AOI22_X1 slo__sro_c2286 (.ZN (slo__sro_n2348), .A1 (n_6_21), .A2 (opt_ipo_n24358)
    , .B1 (n_6_20), .B2 (slo__n30589));
INV_X1 i_6_1_2093 (.ZN (n_6_2907), .A (n_6_1_1106));
AOI22_X1 slo__sro_c2360 (.ZN (slo__sro_n2410), .A1 (n_6_28), .A2 (opt_ipo_n24358)
    , .B1 (drc_ipo_n26574), .B2 (slo__n30589));
INV_X1 i_6_1_2091 (.ZN (n_6_2906), .A (n_6_1_1105));
AOI22_X1 slo__sro_c2247 (.ZN (slo__sro_n2319), .A1 (n_6_22), .A2 (opt_ipo_n24358)
    , .B1 (n_6_21), .B2 (slo__n30589));
INV_X1 i_6_1_2089 (.ZN (n_6_2905), .A (n_6_1_1104));
AOI22_X1 slo__sro_c2147 (.ZN (slo__sro_n2232), .A1 (CLOCK_sgo__n47025), .A2 (opt_ipo_n24358)
    , .B1 (CLOCK_sgo__n47003), .B2 (slo__n30589));
INV_X1 i_6_1_2087 (.ZN (n_6_2904), .A (n_6_1_1103));
AOI22_X1 slo__sro_c2274 (.ZN (slo__sro_n2339), .A1 (n_6_26), .A2 (opt_ipo_n24358)
    , .B1 (n_6_25), .B2 (slo__n30589));
INV_X1 i_6_1_2085 (.ZN (n_6_2903), .A (n_6_1_1102));
AOI21_X4 slo__sro_c38940 (.ZN (slo__sro_n35270), .A (slo__sro_n35271), .B1 (n_6_132), .B2 (n_6_1_1044));
INV_X1 i_6_1_2083 (.ZN (n_6_2902), .A (slo__sro_n2346));
AOI21_X1 slo__sro_c2075 (.ZN (slo__sro_n2166), .A (slo__sro_n2167), .B1 (n_6_12), .B2 (opt_ipo_n24358));
INV_X1 i_6_1_2081 (.ZN (n_6_2901), .A (n_6_1_1100));
NAND2_X1 slo__sro_c2209 (.ZN (slo__sro_n2287), .A1 (slo__n30589), .A2 (n_6_12));
INV_X1 i_6_1_2079 (.ZN (n_6_2900), .A (slo__sro_n2272));
NAND2_X1 slo__sro_c2159 (.ZN (slo__sro_n2244), .A1 (slo__n30589), .A2 (n_6_14));
INV_X1 i_6_1_2077 (.ZN (n_6_2899), .A (slo__sro_n2230));
AOI22_X1 slo__sro_c2185 (.ZN (slo__sro_n2262), .A1 (n_6_16), .A2 (opt_ipo_n24358)
    , .B1 (n_6_15), .B2 (slo__n30589));
INV_X1 i_6_1_2075 (.ZN (n_6_2898), .A (n_6_1_1097));
AOI22_X1 slo__sro_c2197 (.ZN (slo__sro_n2274), .A1 (n_6_19), .A2 (opt_ipo_n24358)
    , .B1 (CLOCK_sgo__n47025), .B2 (slo__n30589));
INV_X1 i_6_1_2073 (.ZN (n_6_2897), .A (slo__sro_n2260));
AOI22_X1 slo__sro_c2173 (.ZN (slo__sro_n2253), .A1 (CLOCK_sgo__n47003), .A2 (opt_ipo_n24358)
    , .B1 (n_6_16), .B2 (slo__n30589));
INV_X1 i_6_1_2071 (.ZN (n_6_2896), .A (n_6_1_1095));
AND2_X1 slo__sro_c2133 (.ZN (slo__sro_n2222), .A1 (n_6_22), .A2 (slo__n30589));
INV_X1 i_6_1_2069 (.ZN (n_6_2895), .A (slo__sro_n2206));
INV_X1 slo__sro_c2231 (.ZN (slo__sro_n2309), .A (CLOCK_sgo__n47054));
INV_X1 i_6_1_2067 (.ZN (n_6_2894), .A (slo__sro_n2284));
AND2_X1 slo__sro_c2119 (.ZN (slo__sro_n2209), .A1 (slo__n30589), .A2 (n_6_13));
INV_X1 i_6_1_2065 (.ZN (n_6_2893), .A (slo__sro_n2164));
AOI21_X1 slo__sro_c2120 (.ZN (slo__sro_n2208), .A (slo__sro_n2209), .B1 (n_6_14), .B2 (opt_ipo_n24358));
INV_X1 i_6_1_2063 (.ZN (n_6_2892), .A (slo__sro_n2194));
AOI22_X1 slo__sro_c2005 (.ZN (slo__sro_n2108), .A1 (n_6_7), .A2 (opt_ipo_n24358), .B1 (drc_ipo_n26594), .B2 (slo__n30589));
INV_X1 i_6_1_2061 (.ZN (n_6_2891), .A (n_6_1_1090));
AND2_X1 slo__sro_c2074 (.ZN (slo__sro_n2167), .A1 (slo__n30589), .A2 (n_6_11));
INV_X1 i_6_1_2059 (.ZN (n_6_2890), .A (n_6_1_1089));
AOI22_X1 sgo__sro_c1500 (.ZN (sgo__sro_n1677), .A1 (n_6_4), .A2 (opt_ipo_n24358), .B1 (n_6_3), .B2 (slo__n30589));
INV_X4 i_6_1_2057 (.ZN (n_6_2889), .A (n_6_1_1088));
AOI22_X1 slo__sro_c2021 (.ZN (slo__sro_n2123), .A1 (n_6_9), .A2 (opt_ipo_n24358), .B1 (n_6_8), .B2 (slo__n30589));
NAND2_X2 CLOCK_slo__sro_c54307 (.ZN (CLOCK_slo__sro_n49673), .A1 (CLOCK_slo__sro_n49674), .A2 (slo__sro_n41144));
INV_X1 sgo__sro_c1550 (.ZN (sgo__sro_n1718), .A (sgo__sro_n1719));
INV_X2 i_6_1_2053 (.ZN (n_6_2887), .A (sgo__sro_n1686));
NAND2_X1 sgo__sro_c1417 (.ZN (sgo__sro_n1602), .A1 (sgo__n711), .A2 (sgo__n1314));
INV_X1 i_6_1_2051 (.ZN (n_6_2886), .A (n_6_1_1085));
AOI22_X1 sgo__sro_c1549 (.ZN (sgo__sro_n1719), .A1 (n_6_10), .A2 (opt_ipo_n24358)
    , .B1 (drc_ipo_n26591), .B2 (slo__n30589));
INV_X1 i_6_1_2049 (.ZN (n_6_2885), .A (slo__sro_n15079));
BUF_X32 slo__c30130 (.Z (slo__n26761), .A (drc_ipo_n26596));
INV_X1 i_6_1_2047 (.ZN (n_6_2884), .A (sgo__sro_n1599));
AOI21_X1 slo__sro_c2051 (.ZN (n_6_1_1100), .A (slo__sro_n2142), .B1 (n_6_51), .B2 (n_6_1_1114));
INV_X2 i_6_1_2045 (.ZN (n_6_2883), .A (sgo__sro_n1557));
AOI22_X1 slo__sro_c2314 (.ZN (slo__sro_n2372), .A1 (drc_ipo_n26574), .A2 (opt_ipo_n24358)
    , .B1 (n_6_26), .B2 (slo__n30589));
NAND2_X1 CLOCK_slo__sro_c53774 (.ZN (CLOCK_slo__sro_n49189), .A1 (CLOCK_slo__sro_n49190), .A2 (CLOCK_slo__sro_n49191));
NOR2_X1 i_6_1_2042 (.ZN (sgo__n675), .A1 (n_6_1_1117), .A2 (Multiplicand[1]));
NOR2_X1 i_6_1_2041 (.ZN (sgo__n687), .A1 (Multiplicand[2]), .A2 (n_6_1_1116));
NOR2_X4 i_6_1_2040 (.ZN (slo__n13799), .A1 (n_6_1_1080), .A2 (n_6_1_1079));
AND2_X1 i_6_1_2039 (.ZN (n_6_1_1077), .A1 (n_6_2912), .A2 (slo__n13799));
AOI221_X1 i_6_1_2038 (.ZN (n_6_1_1076), .A (n_6_1_1077), .B1 (n_6_94), .B2 (n_6_1_1079)
    , .C1 (n_6_126), .C2 (n_6_1_1080));
INV_X1 i_6_1_2037 (.ZN (n_6_2881), .A (n_6_1_1076));
AOI221_X1 i_6_1_2036 (.ZN (n_6_1_1075), .A (n_6_1_1077), .B1 (n_6_93), .B2 (n_6_1_1079)
    , .C1 (n_6_125), .C2 (n_6_1_1080));
INV_X1 i_6_1_2035 (.ZN (n_6_2880), .A (n_6_1_1075));
NAND2_X1 slo__sro_c41188 (.ZN (slo__sro_n37307), .A1 (n_6_1_905), .A2 (n_6_435));
NAND2_X1 slo__sro_c15457 (.ZN (slo__sro_n13955), .A1 (n_6_2648), .A2 (n_6_1_798));
NAND2_X1 slo__sro_c40764 (.ZN (slo__sro_n36945), .A1 (n_6_1_625), .A2 (n_6_932));
NAND2_X1 slo__sro_c5084 (.ZN (slo__sro_n4847), .A1 (n_6_1_238), .A2 (n_6_2160));
INV_X1 i_6_1_2029 (.ZN (n_6_2877), .A (n_6_1_1072));
NAND2_X1 slo__sro_c9054 (.ZN (slo__sro_n8453), .A1 (n_6_2900), .A2 (slo__n13799));
INV_X2 i_6_1_2027 (.ZN (n_6_2876), .A (n_6_1_1071));
NAND2_X1 slo__sro_c8488 (.ZN (slo__sro_n7961), .A1 (n_6_2627), .A2 (n_6_1_763));
INV_X1 i_6_1_2025 (.ZN (n_6_2875), .A (slo__sro_n7944));
NAND2_X1 slo__sro_c8940 (.ZN (slo__sro_n8358), .A1 (slo__n13799), .A2 (n_6_2902));
AOI21_X2 CLOCK_slo__sro_c53775 (.ZN (CLOCK_slo__sro_n49188), .A (CLOCK_slo__sro_n49189)
    , .B1 (n_6_590), .B2 (n_6_1_799));
INV_X1 slo__sro_c23941 (.ZN (slo__sro_n20848), .A (slo__sro_n7448));
INV_X1 i_6_1_2021 (.ZN (n_6_2873), .A (slo__sro_n6519));
AOI222_X2 slo__sro_c8972 (.ZN (slo__sro_n8380), .A1 (n_6_185), .A2 (n_6_1_1045), .B1 (n_6_153)
    , .B2 (n_6_1_1044), .C1 (slo__n18727), .C2 (CLOCK_sgo__n46945));
INV_X1 i_6_1_2019 (.ZN (n_6_2872), .A (n_6_1_1067));
NAND2_X1 slo__sro_c9014 (.ZN (slo__sro_n8417), .A1 (n_6_2901), .A2 (slo__n13799));
INV_X2 i_6_1_2017 (.ZN (n_6_2871), .A (n_6_1_1066));
NAND2_X1 slo__sro_c8956 (.ZN (slo__sro_n8370), .A1 (n_6_2904), .A2 (slo__n13799));
INV_X1 i_6_1_2015 (.ZN (n_6_2870), .A (slo__sro_n39888));
NAND2_X1 slo__sro_c9030 (.ZN (slo__sro_n8432), .A1 (n_6_2908), .A2 (slo__n13799));
INV_X1 i_6_1_2013 (.ZN (n_6_2869), .A (slo__sro_n39898));
AOI222_X1 slo__sro_c9107 (.ZN (slo__sro_n8500), .A1 (n_6_532), .A2 (n_6_1_834), .B1 (n_6_564)
    , .B2 (n_6_1_835), .C1 (n_6_2686), .C2 (CLOCK_sgo__n46922));
INV_X4 i_6_1_2011 (.ZN (n_6_2868), .A (slo__sro_n8450));
AOI21_X2 slo__sro_c33835 (.ZN (slo__sro_n30284), .A (slo__sro_n30285), .B1 (n_6_1131), .B2 (slo___n23268));
INV_X1 i_6_1_2009 (.ZN (n_6_2867), .A (CLOCK_slo__sro_n62530));
INV_X1 i_6_1_2007 (.ZN (n_6_2866), .A (slo__sro_n17238));
INV_X1 slo__sro_c25577 (.ZN (slo__sro_n22350), .A (slo__sro_n15143));
INV_X1 i_6_1_2005 (.ZN (n_6_2865), .A (slo__sro_n22325));
AND2_X1 slo__sro_c24717 (.ZN (slo__sro_n21561), .A1 (n_6_2513), .A2 (n_6_1_658));
INV_X1 i_6_1_2003 (.ZN (n_6_2864), .A (n_6_1_1059));
NOR2_X2 slo__sro_c35873 (.ZN (slo__sro_n32212), .A1 (slo__sro_n32213), .A2 (slo__sro_n10650));
INV_X1 i_6_1_2001 (.ZN (n_6_2863), .A (slo__sro_n32182));
INV_X1 slo__c39499 (.ZN (slo__n35792), .A (n_6_1_1097));
INV_X1 i_6_1_1999 (.ZN (n_6_2862), .A (slo__sro_n35681));
NAND2_X1 CLOCK_slo__sro_c55688 (.ZN (CLOCK_slo__sro_n50913), .A1 (n_6_1258), .A2 (slo___n23274));
INV_X1 i_6_1_1997 (.ZN (n_6_2861), .A (CLOCK_slo__sro_n52568));
AOI221_X2 CLOCK_slo__sro_c58246 (.ZN (slo__sro_n27499), .A (slo__sro_n27500), .B1 (n_6_274)
    , .B2 (n_6_1_974), .C1 (n_6_306), .C2 (n_6_1_975));
INV_X1 i_6_1_1995 (.ZN (n_6_2860), .A (n_6_1_1055));
AOI222_X2 i_6_1_1994 (.ZN (n_6_1_1054), .A1 (n_6_72), .A2 (n_6_1_1079), .B1 (n_6_104)
    , .B2 (n_6_1_1080), .C1 (n_6_2891), .C2 (slo__n13799));
INV_X1 i_6_1_1993 (.ZN (n_6_2859), .A (n_6_1_1054));
AOI21_X2 CLOCK_slo__sro_c59817 (.ZN (slo__sro_n38758), .A (slo__sro_n38759), .B1 (n_6_879), .B2 (n_6_1_660));
INV_X2 i_6_1_1991 (.ZN (n_6_2858), .A (n_6_1_1053));
NAND2_X1 slo__sro_c8998 (.ZN (slo__sro_n8404), .A1 (n_6_2903), .A2 (slo__n13799));
INV_X1 i_6_1_1989 (.ZN (n_6_2857), .A (n_6_1_1052));
NAND2_X1 slo__sro_c9673 (.ZN (slo__sro_n9010), .A1 (slo__n13799), .A2 (n_6_2886));
INV_X2 i_6_1_1987 (.ZN (spw__n68416), .A (slo__sro_n8991));
AOI21_X2 slo__sro_c37896 (.ZN (slo__sro_n34276), .A (slo__sro_n34277), .B1 (n_6_1368), .B2 (n_6_1_379));
INV_X2 i_6_1_1985 (.ZN (n_6_2855), .A (slo__sro_n34136));
AND2_X1 slo__sro_c9758 (.ZN (slo__sro_n9086), .A1 (n_6_2547), .A2 (n_6_1_693));
INV_X4 i_6_1_1983 (.ZN (n_6_2854), .A (slo__sro_n9007));
NAND2_X2 slo__sro_c38939 (.ZN (slo__sro_n35271), .A1 (slo__sro_n35272), .A2 (slo__sro_n8669));
INV_X1 i_6_1_1981 (.ZN (n_6_2853), .A (slo__sro_n8602));
AND2_X1 CLOCK_slo__sro_c64882 (.ZN (CLOCK_slo__sro_n58465), .A1 (n_6_2042), .A2 (n_6_1_98));
INV_X1 i_6_1_1979 (.ZN (n_6_2852), .A (n_6_1_1047));
INV_X2 CLOCK_slo__c59659 (.ZN (CLOCK_slo__n54289), .A (n_6_1_201));
INV_X2 i_6_1_1977 (.ZN (n_6_2851), .A (CLOCK_slo__sro_n61295));
NOR2_X4 i_6_1_1976 (.ZN (sgo__n659), .A1 (n_6_1_1118), .A2 (Multiplicand[2]));
NOR2_X4 i_6_1_1975 (.ZN (sgo__n666), .A1 (Multiplicand[3]), .A2 (n_6_1_1117));
NOR2_X4 i_6_1_1974 (.ZN (CLOCK_sgo__n46945), .A1 (n_6_1_1045), .A2 (n_6_1_1044));
AND2_X1 i_6_1_1973 (.ZN (n_6_1_1042), .A1 (n_6_2881), .A2 (CLOCK_sgo__n46945));
AOI221_X2 i_6_1_1972 (.ZN (n_6_1_1041), .A (n_6_1_1042), .B1 (n_6_190), .B2 (n_6_1_1045)
    , .C1 (n_6_158), .C2 (n_6_1_1044));
INV_X2 i_6_1_1971 (.ZN (n_6_2850), .A (n_6_1_1041));
INV_X2 i_6_1_1969 (.ZN (n_6_2849), .A (n_6_1_1040));
NAND2_X1 slo__sro_c20461 (.ZN (slo__sro_n17953), .A1 (n_6_1_588), .A2 (n_6_2455));
INV_X1 i_6_1_1967 (.ZN (n_6_2848), .A (slo__sro_n40769));
AOI222_X2 i_6_1_1966 (.ZN (n_6_1_1038), .A1 (n_6_187), .A2 (n_6_1_1045), .B1 (n_6_155)
    , .B2 (n_6_1_1044), .C1 (n_6_1_1074), .C2 (CLOCK_sgo__n46945));
INV_X1 i_6_1_1965 (.ZN (n_6_2847), .A (n_6_1_1038));
INV_X2 slo__c39164 (.ZN (slo__n35483), .A (n_6_1_1047));
INV_X2 i_6_1_1963 (.ZN (n_6_2846), .A (n_6_1_1037));
NAND2_X1 slo__sro_c8982 (.ZN (slo__sro_n8392), .A1 (n_6_2889), .A2 (slo__n13799));
INV_X2 i_6_1_1961 (.ZN (n_6_2845), .A (slo__sro_n8380));
NAND2_X1 slo__sro_c35180 (.ZN (slo__sro_n31561), .A1 (n_6_935), .A2 (n_6_1_625));
INV_X1 i_6_1_1959 (.ZN (n_6_2844), .A (n_6_1_1035));
NOR2_X1 slo__sro_c22998 (.ZN (slo__sro_n19971), .A1 (slo__sro_n19973), .A2 (slo__sro_n19972));
INV_X1 i_6_1_1957 (.ZN (n_6_2843), .A (n_6_1_1034));
NAND2_X1 slo__sro_c24342 (.ZN (slo__sro_n21212), .A1 (n_6_2756), .A2 (CLOCK_sgo__n46934));
INV_X1 i_6_1_1955 (.ZN (n_6_2842), .A (CLOCK_slo__sro_n56608));
INV_X1 slo__sro_c11191 (.ZN (slo__sro_n10379), .A (CLOCK_sgo__n46934));
INV_X1 i_6_1_1953 (.ZN (slo___n7881), .A (n_6_1_1032));
AOI21_X2 slo__sro_c33169 (.ZN (slo__sro_n29650), .A (slo__sro_n29651), .B1 (n_6_1317), .B2 (slo___n43257));
INV_X1 i_6_1_1951 (.ZN (n_6_2840), .A (slo__sro_n29523));
NAND2_X1 slo__sro_c41068 (.ZN (slo__sro_n37211), .A1 (n_6_1_763), .A2 (n_6_2629));
INV_X2 i_6_1_1949 (.ZN (n_6_2839), .A (n_6_1_1030));
AOI222_X2 i_6_1_1948 (.ZN (n_6_1_1029), .A1 (n_6_146), .A2 (n_6_1_1044), .B1 (n_6_178)
    , .B2 (n_6_1_1045), .C1 (n_6_2870), .C2 (CLOCK_sgo__n46945));
INV_X2 i_6_1_1947 (.ZN (slo___n8281), .A (n_6_1_1029));
NAND2_X1 slo__sro_c33558 (.ZN (slo__sro_n30034), .A1 (slo__n26894), .A2 (CLOCK_sgo__n46922));
INV_X2 i_6_1_1945 (.ZN (CLOCK_slo___n57806), .A (slo__sro_n29917));
NAND2_X1 slo__sro_c26280 (.ZN (slo__sro_n22965), .A1 (n_6_2213), .A2 (n_6_1_308));
INV_X1 i_6_1_1943 (.ZN (n_6_2836), .A (slo__sro_n37053));
NOR2_X2 slo__sro_c36161 (.ZN (slo__sro_n32484), .A1 (slo__sro_n9873), .A2 (slo__sro_n32485));
INV_X1 i_6_1_1941 (.ZN (n_6_2835), .A (slo__sro_n32357));
NAND2_X2 slo__sro_c33380 (.ZN (slo__sro_n29859), .A1 (n_6_1687), .A2 (n_6_1_204));
INV_X1 i_6_1_1939 (.ZN (n_6_2834), .A (CLOCK_slo__sro_n51306));
NAND2_X1 slo__sro_c24485 (.ZN (slo__sro_n21349), .A1 (n_6_2528), .A2 (n_6_1_658));
INV_X1 i_6_1_1937 (.ZN (n_6_2833), .A (n_6_1_1024));
INV_X1 CLOCK_slo__sro_c54366 (.ZN (CLOCK_slo__sro_n49728), .A (n_6_1_237));
INV_X2 i_6_1_1935 (.ZN (n_6_2832), .A (n_6_1_1023));
AND2_X1 slo__sro_c12819 (.ZN (slo__sro_n11755), .A1 (n_6_2319), .A2 (n_6_1_413));
INV_X1 i_6_1_1933 (.ZN (n_6_2831), .A (slo__sro_n11706));
INV_X1 slo__sro_c24581 (.ZN (slo__sro_n21439), .A (slo__sro_n15779));
INV_X1 i_6_1_1931 (.ZN (n_6_2830), .A (n_6_1_1021));
NAND2_X1 slo__sro_c4982 (.ZN (slo__sro_n4752), .A1 (n_6_1_874), .A2 (n_6_1_868));
INV_X1 i_6_1_1929 (.ZN (n_6_2829), .A (n_6_1_1020));
AOI222_X2 slo__sro_c18228 (.ZN (CLOCK_slo__n50780), .A1 (n_6_243), .A2 (n_6_1_1010)
    , .B1 (n_6_211), .B2 (n_6_1_1009), .C1 (n_6_2840), .C2 (CLOCK_sgo__n46950));
INV_X1 i_6_1_1927 (.ZN (n_6_2828), .A (slo__sro_n16215));
INV_X2 opt_ipo_c27161 (.ZN (opt_ipo_n23778), .A (n_6_1_458));
INV_X2 i_6_1_1925 (.ZN (n_6_2827), .A (n_6_1_1018));
AOI222_X2 i_6_1_1924 (.ZN (n_6_1_1017), .A1 (n_6_134), .A2 (n_6_1_1044), .B1 (n_6_166)
    , .B2 (n_6_1_1045), .C1 (n_6_2858), .C2 (CLOCK_sgo__n46945));
INV_X2 i_6_1_1923 (.ZN (n_6_2826), .A (n_6_1_1017));
INV_X1 CLOCK_slo__sro_c56938 (.ZN (CLOCK_slo__sro_n51982), .A (slo__sro_n5844));
NAND2_X1 CLOCK_slo__sro_c54229 (.ZN (CLOCK_slo__sro_n49603), .A1 (CLOCK_slo__sro_n49604), .A2 (CLOCK_slo__sro_n49605));
NAND2_X1 slo__sro_c9321 (.ZN (slo__sro_n8686), .A1 (n_6_2482), .A2 (n_6_1_623));
NAND2_X1 CLOCK_slo__sro_c54291 (.ZN (CLOCK_slo__sro_n49664), .A1 (n_6_1_378), .A2 (n_6_2271));
NAND2_X1 slo__sro_c10171 (.ZN (slo__sro_n9471), .A1 (n_6_2112), .A2 (n_6_1_203));
NAND2_X4 slo__sro_c33648 (.ZN (slo__sro_n30111), .A1 (slo__sro_n30112), .A2 (slo__sro_n30113));
INV_X1 CLOCK_slo__sro_c55041 (.ZN (CLOCK_slo__sro_n50332), .A (slo__sro_n21561));
INV_X2 i_6_1_1915 (.ZN (slo___n5717), .A (slo__sro_n8949));
NOR2_X1 CLOCK_slo__sro_c57143 (.ZN (CLOCK_slo__sro_n52136), .A1 (slo__sro_n27972), .A2 (CLOCK_slo__sro_n52137));
INV_X2 i_6_1_1913 (.ZN (n_6_2821), .A (CLOCK_slo__sro_n61347));
AOI222_X2 slo__sro_c37381 (.ZN (slo__sro_n33706), .A1 (n_6_756), .A2 (n_6_1_730), .B1 (n_6_724)
    , .B2 (n_6_1_729), .C1 (n_6_2593), .C2 (n_6_1_728));
INV_X2 i_6_1_1911 (.ZN (n_6_2820), .A (slo__sro_n33677));
NOR2_X1 i_6_1_1910 (.ZN (sgo__n644), .A1 (n_6_1_1119), .A2 (Multiplicand[3]));
NOR2_X4 i_6_1_1909 (.ZN (sgo__n656), .A1 (Multiplicand[4]), .A2 (n_6_1_1118));
NOR2_X4 i_6_1_1908 (.ZN (CLOCK_sgo__n46950), .A1 (n_6_1_1010), .A2 (n_6_1_1009));
AND2_X1 i_6_1_1907 (.ZN (n_6_1_1007), .A1 (n_6_2850), .A2 (CLOCK_sgo__n46950));
AOI221_X2 i_6_1_1906 (.ZN (n_6_1_1006), .A (n_6_1_1007), .B1 (n_6_222), .B2 (n_6_1_1009)
    , .C1 (n_6_254), .C2 (n_6_1_1010));
AOI21_X2 CLOCK_sgo__sro_c51594 (.ZN (slo__sro_n5416), .A (CLOCK_sgo__sro_n47337), .B1 (n_6_582), .B2 (n_6_1_799));
NAND2_X1 slo__sro_c26010 (.ZN (slo__sro_n22736), .A1 (n_6_2780), .A2 (CLOCK_sgo__n46937));
INV_X4 i_6_1_1903 (.ZN (n_6_2818), .A (slo__sro_n22701));
NAND2_X1 slo__sro_c12635 (.ZN (slo__sro_n11597), .A1 (n_6_2322), .A2 (n_6_1_413));
INV_X1 i_6_1_1901 (.ZN (n_6_2817), .A (n_6_1_1004));
INV_X1 i_6_1_1899 (.ZN (n_6_2816), .A (slo__sro_n41830));
AND2_X1 slo__sro_c12913 (.ZN (slo__sro_n11844), .A1 (n_6_2349), .A2 (n_6_1_448));
INV_X2 i_6_1_1897 (.ZN (n_6_2815), .A (slo__sro_n20612));
NAND2_X1 slo__sro_c25976 (.ZN (slo__sro_n22703), .A1 (n_6_253), .A2 (n_6_1_1010));
INV_X1 i_6_1_1895 (.ZN (slo___n18581), .A (n_6_1_1001));
NAND2_X1 slo__sro_c34812 (.ZN (slo__sro_n31219), .A1 (slo___n23364), .A2 (n_6_1180));
INV_X2 i_6_1_1893 (.ZN (n_6_2813), .A (n_6_1_1000));
NAND2_X1 slo__sro_c41383 (.ZN (slo__sro_n37485), .A1 (n_6_2711), .A2 (n_6_1_868));
INV_X1 i_6_1_1891 (.ZN (n_6_2812), .A (slo__sro_n11578));
NAND2_X1 CLOCK_slo__sro_c55257 (.ZN (CLOCK_slo__sro_n50525), .A1 (n_6_1_483), .A2 (n_6_2366));
INV_X2 i_6_1_1889 (.ZN (n_6_2811), .A (n_6_1_998));
NAND2_X1 slo__sro_c24793 (.ZN (slo__sro_n21633), .A1 (n_6_818), .A2 (n_6_1_695));
INV_X1 i_6_1_1887 (.ZN (n_6_2810), .A (slo__sro_n13965));
INV_X1 slo__c18115 (.ZN (slo__n16143), .A (slo__sro_n6762));
INV_X2 i_6_1_1885 (.ZN (n_6_2809), .A (CLOCK_slo__sro_n56057));
NAND2_X1 slo__sro_c18238 (.ZN (slo__sro_n16242), .A1 (n_6_2644), .A2 (n_6_1_798));
NAND2_X1 CLOCK_slo__sro_c55542 (.ZN (CLOCK_slo__sro_n50794), .A1 (n_6_2842), .A2 (CLOCK_sgo__n46950));
NAND2_X1 CLOCK_slo__sro_c62145 (.ZN (CLOCK_slo__sro_n56379), .A1 (n_6_2688), .A2 (CLOCK_sgo__n46922));
INV_X2 i_6_1_1881 (.ZN (n_6_2807), .A (n_6_1_994));
NOR2_X4 CLOCK_slo__sro_c63354 (.ZN (n_6_1_164), .A1 (slo__sro_n13370), .A2 (CLOCK_slo__sro_n57315));
OAI21_X1 slo__mro_c36884 (.ZN (slo__mro_n33237), .A (slo__sro_n20509), .B1 (slo__mro_n33239), .B2 (slo__mro_n33238));
AOI222_X2 i_6_1_1878 (.ZN (n_6_1_992), .A1 (n_6_208), .A2 (n_6_1_1009), .B1 (n_6_240)
    , .B2 (n_6_1_1010), .C1 (CLOCK_slo___n57806), .C2 (CLOCK_sgo__n46950));
INV_X2 i_6_1_1877 (.ZN (n_6_2805), .A (n_6_1_992));
AOI222_X2 i_6_1_1876 (.ZN (n_6_1_991), .A1 (n_6_207), .A2 (n_6_1_1009), .B1 (n_6_239)
    , .B2 (n_6_1_1010), .C1 (n_6_2836), .C2 (CLOCK_sgo__n46950));
INV_X2 i_6_1_1875 (.ZN (n_6_2804), .A (n_6_1_991));
NAND2_X1 CLOCK_slo__sro_c65795 (.ZN (CLOCK_slo__sro_n59304), .A1 (n_6_2306), .A2 (n_6_1_413));
INV_X1 i_6_1_1873 (.ZN (n_6_2803), .A (CLOCK_slo__sro_n59280));
AOI21_X1 CLOCK_slo__sro_c69382 (.ZN (CLOCK_slo__sro_n62488), .A (CLOCK_slo__sro_n49216)
    , .B1 (n_6_490), .B2 (n_6_1_870));
INV_X1 i_6_1_1871 (.ZN (n_6_2802), .A (CLOCK_slo__sro_n62128));
NAND2_X1 slo__sro_c21048 (.ZN (slo__sro_n18405), .A1 (slo___n23215), .A2 (n_6_1614));
INV_X1 i_6_1_1869 (.ZN (n_6_2801), .A (CLOCK_slo__sro_n65088));
AOI21_X4 slo__sro_c39193 (.ZN (slo__sro_n35509), .A (slo__sro_n8603), .B1 (n_6_66), .B2 (n_6_1_1079));
INV_X1 i_6_1_1867 (.ZN (n_6_2800), .A (slo__sro_n35466));
NAND2_X1 slo__sro_c35680 (.ZN (slo__sro_n32027), .A1 (slo__sro_n32029), .A2 (slo__sro_n32028));
INV_X2 i_6_1_1865 (.ZN (n_6_2799), .A (slo__sro_n31830));
NAND2_X1 slo__sro_c9301 (.ZN (slo__sro_n8669), .A1 (n_6_2856), .A2 (CLOCK_sgo__n46945));
NAND2_X1 CLOCK_sgo__sro_c52079 (.ZN (CLOCK_sgo__sro_n47734), .A1 (n_6_1_308), .A2 (n_6_2206));
AOI222_X2 i_6_1_1862 (.ZN (CLOCK_slo__n62554), .A1 (n_6_200), .A2 (n_6_1_1009), .B1 (n_6_232)
    , .B2 (n_6_1_1010), .C1 (n_6_2829), .C2 (CLOCK_sgo__n46950));
NAND2_X1 CLOCK_slo__sro_c69578 (.ZN (CLOCK_slo__sro_n62669), .A1 (opt_ipo_n24285), .A2 (n_6_1_658));
AOI222_X2 i_6_1_1860 (.ZN (n_6_1_983), .A1 (n_6_199), .A2 (n_6_1_1009), .B1 (n_6_231)
    , .B2 (n_6_1_1010), .C1 (n_6_2828), .C2 (CLOCK_sgo__n46950));
INV_X2 i_6_1_1859 (.ZN (n_6_2796), .A (n_6_1_983));
NAND2_X1 CLOCK_slo__sro_c68486 (.ZN (CLOCK_slo__sro_n61697), .A1 (n_6_1_1079), .A2 (n_6_68));
INV_X2 i_6_1_1857 (.ZN (n_6_2795), .A (slo__sro_n35197));
INV_X1 slo__sro_c37456 (.ZN (slo__sro_n33777), .A (slo__sro_n33778));
INV_X2 i_6_1_1855 (.ZN (n_6_2794), .A (slo__sro_n33755));
NAND2_X1 slo__sro_c8351 (.ZN (slo__sro_n7835), .A1 (n_6_2910), .A2 (slo__n13799));
INV_X2 i_6_1_1853 (.ZN (n_6_2793), .A (slo__sro_n7772));
NAND2_X1 slo__sro_c13155 (.ZN (slo__sro_n12060), .A1 (n_6_2632), .A2 (n_6_1_763));
INV_X2 i_6_1_1851 (.ZN (n_6_2792), .A (n_6_1_979));
AND2_X1 slo__sro_c23741 (.ZN (slo__sro_n20666), .A1 (n_6_2167), .A2 (n_6_1_238));
INV_X1 i_6_1_1849 (.ZN (n_6_2791), .A (slo__sro_n11796));
INV_X2 CLOCK_slo__c62028 (.ZN (CLOCK_slo__n56284), .A (CLOCK_slo__sro_n55447));
INV_X2 i_6_1_1847 (.ZN (n_6_2790), .A (CLOCK_slo__sro_n65030));
AOI221_X2 CLOCK_slo__sro_c64865 (.ZN (n_6_1_1047), .A (CLOCK_slo__sro_n58451), .B1 (n_6_97)
    , .B2 (n_6_1_1080), .C1 (n_6_65), .C2 (n_6_1_1079));
INV_X1 i_6_1_1845 (.ZN (CLOCK_slo___n65042), .A (n_6_1_976));
NOR2_X4 i_6_1_1844 (.ZN (sgo__n630), .A1 (n_6_1_1120), .A2 (Multiplicand[4]));
NOR2_X4 i_6_1_1843 (.ZN (sgo__n637), .A1 (Multiplicand[5]), .A2 (n_6_1_1119));
NOR2_X1 i_6_1_1842 (.ZN (CLOCK_sgo__n46942), .A1 (n_6_1_975), .A2 (n_6_1_974));
AND2_X1 i_6_1_1841 (.ZN (n_6_1_972), .A1 (opt_ipo_n25006), .A2 (n_6_1_973));
AOI221_X2 i_6_1_1840 (.ZN (n_6_1_971), .A (n_6_1_972), .B1 (n_6_286), .B2 (n_6_1_974)
    , .C1 (n_6_318), .C2 (n_6_1_975));
INV_X1 i_6_1_1839 (.ZN (n_6_2788), .A (n_6_1_971));
AOI221_X2 i_6_1_1838 (.ZN (n_6_1_970), .A (n_6_1_972), .B1 (n_6_285), .B2 (n_6_1_974)
    , .C1 (n_6_317), .C2 (n_6_1_975));
INV_X2 i_6_1_1837 (.ZN (n_6_2787), .A (n_6_1_970));
BUF_X32 slo__c35338 (.Z (slo__n31700), .A (drc_ipo_n26597));
INV_X1 i_6_1_1835 (.ZN (n_6_2786), .A (n_6_1_969));
AOI222_X2 i_6_1_1834 (.ZN (n_6_1_968), .A1 (n_6_315), .A2 (n_6_1_975), .B1 (n_6_283)
    , .B2 (n_6_1_974), .C1 (n_6_2817), .C2 (n_6_1_973));
INV_X1 i_6_1_1833 (.ZN (n_6_2785), .A (n_6_1_968));
NAND2_X1 slo__sro_c22403 (.ZN (slo__sro_n19423), .A1 (n_6_2314), .A2 (n_6_1_413));
INV_X1 i_6_1_1831 (.ZN (n_6_2784), .A (n_6_1_967));
BUF_X16 slo__c21753 (.Z (slo__n18930), .A (sgo__n1292));
NAND2_X1 CLOCK_slo__sro_c54368 (.ZN (CLOCK_slo__sro_n49726), .A1 (CLOCK_slo__sro_n49727), .A2 (CLOCK_slo__sro_n49728));
AOI21_X4 slo__sro_c12868 (.ZN (slo__sro_n11796), .A (slo__sro_n11797), .B1 (n_6_194), .B2 (n_6_1_1009));
INV_X2 i_6_1_1827 (.ZN (n_6_2782), .A (n_6_1_965));
INV_X1 slo__c16789 (.ZN (slo__n15087), .A (slo__sro_n11578));
INV_X2 i_6_1_1825 (.ZN (n_6_2781), .A (CLOCK_slo__sro_n53339));
AND2_X1 slo__sro_c17486 (.ZN (slo__sro_n15657), .A1 (slo__sro_n2968), .A2 (n_6_1_308));
INV_X2 i_6_1_1823 (.ZN (n_6_2780), .A (slo__sro_n15586));
AOI222_X2 i_6_1_1822 (.ZN (n_6_1_962), .A1 (n_6_277), .A2 (n_6_1_974), .B1 (n_6_309)
    , .B2 (n_6_1_975), .C1 (n_6_2811), .C2 (n_6_1_973));
INV_X2 i_6_1_1821 (.ZN (n_6_2779), .A (n_6_1_962));
AOI21_X4 slo__sro_c39309 (.ZN (n_6_1_909), .A (slo__sro_n35616), .B1 (n_6_323), .B2 (n_6_1_939));
INV_X1 i_6_1_1819 (.ZN (n_6_2778), .A (slo__sro_n35288));
BUF_X32 drc_ipo_c29975 (.Z (drc_ipo_n26598), .A (slo__n18930));
INV_X1 i_6_1_1817 (.ZN (n_6_2777), .A (n_6_1_960));
NAND2_X1 slo__sro_c30990 (.ZN (slo__sro_n27583), .A1 (n_6_729), .A2 (n_6_1_729));
INV_X2 i_6_1_1815 (.ZN (n_6_2776), .A (slo__sro_n27499));
AOI21_X1 slo__sro_c25143 (.ZN (slo__sro_n21941), .A (slo__sro_n12963), .B1 (n_6_597), .B2 (n_6_1_799));
INV_X1 i_6_1_1813 (.ZN (n_6_2775), .A (CLOCK_slo__sro_n59027));
NAND2_X1 slo__sro_c10236 (.ZN (slo__sro_n9535), .A1 (n_6_1_378), .A2 (n_6_2289));
INV_X2 i_6_1_1811 (.ZN (n_6_2774), .A (slo__sro_n22431));
AOI221_X2 slo__sro_c12504 (.ZN (n_6_1_891), .A (slo__sro_n11483), .B1 (n_6_404), .B2 (n_6_1_904)
    , .C1 (n_6_436), .C2 (n_6_1_905));
INV_X1 i_6_1_1809 (.ZN (n_6_2773), .A (n_6_1_956));
NAND2_X1 slo__sro_c11068 (.ZN (slo__sro_n10271), .A1 (slo__sro_n10272), .A2 (slo__sro_n10273));
INV_X1 i_6_1_1807 (.ZN (n_6_2772), .A (slo__sro_n29674));
INV_X1 slo__c11965 (.ZN (slo__n11048), .A (n_6_1_802));
INV_X1 i_6_1_1805 (.ZN (n_6_2771), .A (slo__sro_n11034));
NAND2_X1 slo__sro_c11987 (.ZN (slo__sro_n11071), .A1 (CLOCK_opt_ipo_n46124), .A2 (n_6_1_868));
INV_X1 i_6_1_1803 (.ZN (n_6_2770), .A (CLOCK_slo__sro_n50068));
AND2_X1 slo__sro_c12001 (.ZN (slo__sro_n11080), .A1 (slo__sro_n34940), .A2 (CLOCK_sgo__n46937));
INV_X1 i_6_1_1801 (.ZN (n_6_2769), .A (slo__sro_n10838));
NAND2_X1 slo__sro_c10431 (.ZN (slo__sro_n9713), .A1 (n_6_2794), .A2 (n_6_1_973));
INV_X1 i_6_1_1799 (.ZN (n_6_2768), .A (n_6_1_951));
NAND2_X1 slo__sro_c26502 (.ZN (slo__sro_n23160), .A1 (n_6_91), .A2 (n_6_1_1079));
INV_X1 i_6_1_1797 (.ZN (n_6_2767), .A (n_6_1_950));
NAND2_X1 slo__sro_c9194 (.ZN (slo__sro_n8582), .A1 (n_6_2899), .A2 (slo__n13799));
INV_X1 i_6_1_1795 (.ZN (n_6_2766), .A (n_6_1_949));
NAND2_X1 slo__sro_c9566 (.ZN (slo__sro_n8903), .A1 (n_6_2371), .A2 (n_6_1_483));
NAND2_X1 CLOCK_slo__sro_c62435 (.ZN (CLOCK_slo__sro_n56598), .A1 (CLOCK_sgo__n46922), .A2 (n_6_2692));
INV_X1 slo__sro_c38854 (.ZN (slo__sro_n35198), .A (slo__sro_n35199));
INV_X2 CLOCK_slo__c53120 (.ZN (slo__sro_n6239), .A (CLOCK_slo__n48618));
INV_X1 CLOCK_slo__sro_c69871 (.ZN (CLOCK_slo__sro_n62932), .A (slo__sro_n19728));
INV_X1 i_6_1_1789 (.ZN (n_6_2763), .A (n_6_1_946));
AOI222_X2 slo__sro_c10542 (.ZN (slo__sro_n9805), .A1 (n_6_1169), .A2 (slo___n23364)
    , .B1 (n_6_1201), .B2 (slo___n23466), .C1 (CLOCK_slo__n55511), .C2 (n_6_1_483));
INV_X1 i_6_1_1787 (.ZN (n_6_2762), .A (n_6_1_945));
NAND2_X1 slo__sro_c31275 (.ZN (slo__sro_n27862), .A1 (n_6_2613), .A2 (n_6_1_763));
NAND2_X1 slo__sro_c35273 (.ZN (slo__sro_n31645), .A1 (n_6_281), .A2 (n_6_1_974));
AOI21_X2 CLOCK_slo__sro_c57131 (.ZN (CLOCK_slo__sro_n52124), .A (CLOCK_slo__sro_n52125)
    , .B1 (n_6_1213), .B2 (slo___n23466));
INV_X4 i_6_1_1783 (.ZN (n_6_2760), .A (n_6_1_943));
AOI222_X2 i_6_1_1782 (.ZN (n_6_1_942), .A1 (n_6_257), .A2 (n_6_1_974), .B1 (n_6_289)
    , .B2 (n_6_1_975), .C1 (n_6_2791), .C2 (n_6_1_973));
INV_X2 i_6_1_1781 (.ZN (CLOCK_slo___n58400), .A (n_6_1_942));
AOI222_X1 i_6_1_1780 (.ZN (n_6_1_941), .A1 (n_6_256), .A2 (n_6_1_974), .B1 (n_6_288)
    , .B2 (n_6_1_975), .C1 (n_6_2790), .C2 (n_6_1_973));
INV_X1 i_6_1_1779 (.ZN (n_6_2758), .A (n_6_1_941));
NOR2_X4 i_6_1_1778 (.ZN (sgo__n618), .A1 (n_6_1_1121), .A2 (Multiplicand[5]));
NOR2_X4 i_6_1_1777 (.ZN (sgo__n621), .A1 (Multiplicand[6]), .A2 (n_6_1_1120));
NOR2_X4 i_6_1_1776 (.ZN (CLOCK_sgo__n46937), .A1 (n_6_1_940), .A2 (n_6_1_939));
AND2_X1 i_6_1_1775 (.ZN (n_6_1_937), .A1 (n_6_2788), .A2 (CLOCK_sgo__n46937));
AOI221_X1 i_6_1_1774 (.ZN (n_6_1_936), .A (n_6_1_937), .B1 (n_6_350), .B2 (n_6_1_939)
    , .C1 (n_6_382), .C2 (n_6_1_940));
INV_X1 i_6_1_1773 (.ZN (n_6_2757), .A (n_6_1_936));
AOI221_X1 i_6_1_1772 (.ZN (n_6_1_935), .A (n_6_1_937), .B1 (n_6_349), .B2 (n_6_1_939)
    , .C1 (n_6_381), .C2 (n_6_1_940));
INV_X1 i_6_1_1771 (.ZN (n_6_2756), .A (n_6_1_935));
NAND2_X1 CLOCK_slo__sro_c66263 (.ZN (CLOCK_slo__sro_n59729), .A1 (n_6_1_100), .A2 (n_6_1911));
INV_X2 i_6_1_1769 (.ZN (n_6_2755), .A (CLOCK_slo__sro_n59712));
AOI222_X2 i_6_1_1768 (.ZN (n_6_1_933), .A1 (n_6_379), .A2 (n_6_1_940), .B1 (n_6_347)
    , .B2 (n_6_1_939), .C1 (n_6_2786), .C2 (CLOCK_sgo__n46937));
INV_X2 i_6_1_1767 (.ZN (n_6_2754), .A (n_6_1_933));
NAND2_X1 slo__sro_c9657 (.ZN (slo__sro_n8994), .A1 (slo__n13799), .A2 (CLOCK_opt_ipo_n46146));
INV_X2 opt_ipo_c49667 (.ZN (opt_ipo_n45324), .A (slo__sro_n6479));
AOI222_X2 i_6_1_1764 (.ZN (n_6_1_931), .A1 (n_6_377), .A2 (n_6_1_940), .B1 (n_6_345)
    , .B2 (n_6_1_939), .C1 (n_6_2784), .C2 (CLOCK_sgo__n46937));
INV_X1 i_6_1_1763 (.ZN (n_6_2752), .A (n_6_1_931));
NAND2_X1 slo__sro_c31398 (.ZN (slo__sro_n27972), .A1 (slo__sro_n27973), .A2 (slo__sro_n27974));
INV_X2 i_6_1_1761 (.ZN (n_6_2751), .A (n_6_1_930));
AND2_X1 slo__sro_c23119 (.ZN (slo__sro_n20081), .A1 (n_6_2134), .A2 (n_6_1_203));
INV_X1 i_6_1_1759 (.ZN (n_6_2750), .A (n_6_1_929));
NAND2_X1 CLOCK_slo__sro_c53148 (.ZN (CLOCK_slo__sro_n48636), .A1 (n_6_485), .A2 (n_6_1_870));
INV_X1 i_6_1_1757 (.ZN (n_6_2749), .A (slo__sro_n11828));
NAND2_X1 slo__sro_c26022 (.ZN (slo__sro_n22745), .A1 (n_6_2530), .A2 (n_6_1_658));
INV_X2 i_6_1_1755 (.ZN (n_6_2748), .A (n_6_1_927));
NAND2_X1 slo__sro_c12866 (.ZN (slo__sro_n11798), .A1 (n_6_226), .A2 (n_6_1_1010));
INV_X1 i_6_1_1753 (.ZN (n_6_2747), .A (n_6_1_926));
INV_X1 slo__sro_c26075 (.ZN (slo__sro_n22780), .A (n_6_1_974));
INV_X1 i_6_1_1751 (.ZN (n_6_2746), .A (n_6_1_925));
NAND2_X1 CLOCK_slo__sro_c54051 (.ZN (CLOCK_slo__sro_n49429), .A1 (n_6_2713), .A2 (n_6_1_868));
INV_X1 i_6_1_1749 (.ZN (n_6_2745), .A (slo__sro_n27391));
INV_X2 slo__c12415 (.ZN (slo__n11409), .A (n_6_1_1001));
INV_X1 i_6_1_1747 (.ZN (n_6_2744), .A (n_6_1_923));
AOI21_X1 slo__sro_c25977 (.ZN (slo__sro_n22702), .A (n_6_1_1007), .B1 (n_6_221), .B2 (n_6_1_1009));
INV_X1 i_6_1_1745 (.ZN (n_6_2743), .A (slo__sro_n22677));
AND2_X1 slo__sro_c5697 (.ZN (slo__sro_n5417), .A1 (n_6_2641), .A2 (n_6_1_798));
INV_X1 i_6_1_1743 (.ZN (n_6_2742), .A (CLOCK_slo__sro_n59773));
INV_X1 slo__c17183 (.ZN (slo__n15402), .A (n_6_1_148));
INV_X1 i_6_1_1741 (.ZN (n_6_2741), .A (n_6_1_920));
INV_X4 CLOCK_slo__c63346 (.ZN (CLOCK_slo__n57308), .A (slo__sro_n19627));
INV_X1 i_6_1_1739 (.ZN (n_6_2740), .A (n_6_1_919));
AOI222_X2 slo__sro_c13485 (.ZN (n_6_1_877), .A1 (n_6_422), .A2 (n_6_1_905), .B1 (n_6_390)
    , .B2 (n_6_1_904), .C1 (opt_ipo_n25116), .C2 (CLOCK_sgo__n46934));
INV_X1 i_6_1_1737 (.ZN (n_6_2739), .A (CLOCK_slo__sro_n51957));
AND2_X1 slo__sro_c23193 (.ZN (slo__sro_n20147), .A1 (n_6_2270), .A2 (n_6_1_378));
INV_X2 i_6_1_1735 (.ZN (n_6_2738), .A (n_6_1_917));
AND2_X1 slo__sro_c10120 (.ZN (slo__sro_n9421), .A1 (n_6_2040), .A2 (n_6_1_98));
INV_X1 i_6_1_1733 (.ZN (n_6_2737), .A (slo__sro_n9341));
AOI221_X2 slo__sro_c9759 (.ZN (slo__sro_n9085), .A (slo__sro_n9086), .B1 (n_6_805)
    , .B2 (n_6_1_695), .C1 (n_6_773), .C2 (n_6_1_694));
INV_X1 i_6_1_1731 (.ZN (n_6_2736), .A (n_6_1_915));
NAND2_X1 slo__sro_c16899 (.ZN (slo__sro_n15183), .A1 (slo__sro_n15184), .A2 (slo__sro_n15185));
INV_X4 i_6_1_1729 (.ZN (n_6_2735), .A (slo__sro_n22347));
NAND2_X1 slo__sro_c8920 (.ZN (slo__sro_n8338), .A1 (slo__sro_n8339), .A2 (slo__sro_n8340));
INV_X1 slo__c16184 (.ZN (slo__n14568), .A (slo__sro_n28562));
NAND2_X1 CLOCK_sgo__sro_c51863 (.ZN (CLOCK_sgo__sro_n47560), .A1 (CLOCK_sgo__sro_n47561), .A2 (CLOCK_sgo__sro_n47562));
NAND2_X1 slo__sro_c12062 (.ZN (slo__sro_n11126), .A1 (n_6_2361), .A2 (n_6_1_483));
INV_X2 i_6_1_1723 (.ZN (n_6_2732), .A (n_6_1_911));
NAND2_X1 slo__sro_c8473 (.ZN (slo__sro_n7946), .A1 (n_6_1_1080), .A2 (n_6_120));
INV_X4 i_6_1_1721 (.ZN (n_6_2731), .A (CLOCK_sgo__sro_n47197));
AND2_X1 slo__sro_c8739 (.ZN (slo__sro_n8180), .A1 (n_6_2475), .A2 (n_6_1_588));
INV_X1 i_6_1_1719 (.ZN (n_6_2730), .A (n_6_1_909));
BUF_X32 drc_ipo_c29960 (.Z (drc_ipo_n26583), .A (CLOCK_sgo__n47002));
INV_X1 i_6_1_1717 (.ZN (n_6_2729), .A (slo__sro_n32138));
AOI222_X1 i_6_1_1716 (.ZN (n_6_1_907), .A1 (n_6_321), .A2 (n_6_1_939), .B1 (n_6_353)
    , .B2 (n_6_1_940), .C1 (n_6_2760), .C2 (CLOCK_sgo__n46937));
INV_X1 i_6_1_1715 (.ZN (n_6_2728), .A (n_6_1_907));
AOI221_X2 slo__sro_c42823 (.ZN (slo__sro_n38698), .A (slo__sro_n38699), .B1 (n_6_1178)
    , .B2 (slo___n23364), .C1 (n_6_1210), .C2 (slo___n23466));
INV_X2 i_6_1_1713 (.ZN (n_6_2727), .A (n_6_1_906));
NOR2_X4 i_6_1_1712 (.ZN (sgo__n610), .A1 (n_6_1_1122), .A2 (Multiplicand[6]));
NOR2_X4 i_6_1_1711 (.ZN (sgo__n613), .A1 (Multiplicand[7]), .A2 (n_6_1_1121));
NOR2_X4 i_6_1_1710 (.ZN (CLOCK_sgo__n46934), .A1 (n_6_1_905), .A2 (n_6_1_904));
AND2_X1 i_6_1_1709 (.ZN (n_6_1_902), .A1 (n_6_2757), .A2 (CLOCK_sgo__n46934));
AOI221_X1 i_6_1_1708 (.ZN (n_6_1_901), .A (n_6_1_902), .B1 (n_6_414), .B2 (n_6_1_904)
    , .C1 (n_6_446), .C2 (n_6_1_905));
INV_X1 i_6_1_1707 (.ZN (n_6_2726), .A (n_6_1_901));
AOI221_X1 i_6_1_1706 (.ZN (n_6_1_900), .A (n_6_1_902), .B1 (n_6_413), .B2 (n_6_1_904)
    , .C1 (n_6_445), .C2 (n_6_1_905));
INV_X1 i_6_1_1705 (.ZN (n_6_2725), .A (n_6_1_900));
NAND2_X1 slo__sro_c24452 (.ZN (slo__sro_n21317), .A1 (n_6_2752), .A2 (CLOCK_sgo__n46934));
INV_X4 i_6_1_1703 (.ZN (n_6_2724), .A (slo__sro_n30704));
NAND2_X1 slo__sro_c11529 (.ZN (slo__sro_n10650), .A1 (slo__sro_n10651), .A2 (slo__sro_n10652));
INV_X4 i_6_1_1701 (.ZN (n_6_2723), .A (n_6_1_898));
NAND2_X1 slo__sro_c33559 (.ZN (slo__sro_n30033), .A1 (n_6_1_835), .A2 (n_6_565));
INV_X1 i_6_1_1699 (.ZN (n_6_2722), .A (slo__sro_n34606));
INV_X1 slo__sro_c9644 (.ZN (slo__sro_n8978), .A (slo__sro_n8979));
INV_X4 i_6_1_1697 (.ZN (n_6_2721), .A (slo__sro_n8965));
AND2_X1 slo__sro_c9496 (.ZN (slo__sro_n8834), .A1 (n_6_2600), .A2 (n_6_1_728));
INV_X1 i_6_1_1695 (.ZN (n_6_2720), .A (slo__sro_n21314));
NAND2_X1 slo__sro_c11257 (.ZN (slo__sro_n10427), .A1 (slo__sro_n10428), .A2 (slo__sro_n10429));
INV_X1 i_6_1_1693 (.ZN (n_6_2719), .A (n_6_1_894));
AOI222_X2 slo__sro_c8086 (.ZN (n_6_1_815), .A1 (n_6_558), .A2 (n_6_1_835), .B1 (n_6_526)
    , .B2 (n_6_1_834), .C1 (n_6_2680), .C2 (CLOCK_sgo__n46922));
INV_X1 i_6_1_1691 (.ZN (n_6_2718), .A (slo__sro_n7583));
AOI222_X2 i_6_1_1690 (.ZN (n_6_1_892), .A1 (n_6_437), .A2 (n_6_1_905), .B1 (n_6_405)
    , .B2 (n_6_1_904), .C1 (n_6_2749), .C2 (CLOCK_sgo__n46934));
INV_X2 i_6_1_1689 (.ZN (n_6_2717), .A (n_6_1_892));
AOI222_X1 slo__sro_c12523 (.ZN (slo__sro_n11496), .A1 (n_6_1862), .A2 (n_6_1_99), .B1 (n_6_1894)
    , .B2 (n_6_1_100), .C1 (n_6_2021), .C2 (n_6_1_98));
INV_X2 i_6_1_1687 (.ZN (n_6_2716), .A (n_6_1_891));
AND2_X1 CLOCK_slo__sro_c56461 (.ZN (CLOCK_slo__sro_n51595), .A1 (n_6_2088), .A2 (n_6_1_168));
INV_X2 i_6_1_1685 (.ZN (n_6_2715), .A (CLOCK_slo__sro_n60125));
INV_X1 slo__c15442 (.ZN (slo__n13938), .A (slo__sro_n9075));
INV_X2 i_6_1_1683 (.ZN (n_6_2714), .A (slo__sro_n35375));
NAND2_X1 slo__sro_c33443 (.ZN (slo__sro_n29919), .A1 (n_6_2869), .A2 (CLOCK_sgo__n46945));
INV_X2 i_6_1_1681 (.ZN (n_6_2713), .A (n_6_1_888));
AOI222_X2 i_6_1_1680 (.ZN (n_6_1_887), .A1 (n_6_400), .A2 (n_6_1_904), .B1 (n_6_432)
    , .B2 (n_6_1_905), .C1 (n_6_2744), .C2 (CLOCK_sgo__n46934));
INV_X1 i_6_1_1679 (.ZN (n_6_2712), .A (n_6_1_887));
AOI222_X2 i_6_1_1678 (.ZN (n_6_1_886), .A1 (n_6_399), .A2 (n_6_1_904), .B1 (n_6_431)
    , .B2 (n_6_1_905), .C1 (n_6_2743), .C2 (CLOCK_sgo__n46934));
INV_X2 i_6_1_1677 (.ZN (n_6_2711), .A (n_6_1_886));
AOI222_X1 i_6_1_1676 (.ZN (n_6_1_885), .A1 (n_6_398), .A2 (n_6_1_904), .B1 (n_6_430)
    , .B2 (n_6_1_905), .C1 (n_6_2742), .C2 (CLOCK_sgo__n46934));
INV_X1 i_6_1_1675 (.ZN (n_6_2710), .A (n_6_1_885));
AOI222_X2 i_6_1_1674 (.ZN (n_6_1_884), .A1 (n_6_397), .A2 (n_6_1_904), .B1 (n_6_429)
    , .B2 (n_6_1_905), .C1 (n_6_2741), .C2 (CLOCK_sgo__n46934));
INV_X1 i_6_1_1673 (.ZN (n_6_2709), .A (n_6_1_884));
AOI222_X1 i_6_1_1672 (.ZN (n_6_1_883), .A1 (n_6_396), .A2 (n_6_1_904), .B1 (n_6_428)
    , .B2 (n_6_1_905), .C1 (n_6_2740), .C2 (CLOCK_sgo__n46934));
INV_X1 i_6_1_1671 (.ZN (slo___n16308), .A (n_6_1_883));
AOI222_X1 i_6_1_1670 (.ZN (n_6_1_882), .A1 (n_6_395), .A2 (n_6_1_904), .B1 (n_6_427)
    , .B2 (n_6_1_905), .C1 (n_6_2739), .C2 (CLOCK_sgo__n46934));
INV_X1 i_6_1_1669 (.ZN (n_6_2707), .A (n_6_1_882));
AOI222_X1 i_6_1_1668 (.ZN (n_6_1_881), .A1 (n_6_394), .A2 (n_6_1_904), .B1 (n_6_426)
    , .B2 (n_6_1_905), .C1 (n_6_2738), .C2 (CLOCK_sgo__n46934));
INV_X1 i_6_1_1667 (.ZN (slo___n8747), .A (n_6_1_881));
AOI222_X2 i_6_1_1666 (.ZN (n_6_1_880), .A1 (n_6_393), .A2 (n_6_1_904), .B1 (n_6_425)
    , .B2 (n_6_1_905), .C1 (n_6_2737), .C2 (CLOCK_sgo__n46934));
AOI221_X2 slo__sro_c33445 (.ZN (slo__sro_n29917), .A (slo__sro_n29918), .B1 (n_6_177)
    , .B2 (n_6_1_1045), .C1 (n_6_145), .C2 (n_6_1_1044));
BUF_X2 CLOCK_slo___L1_c72228 (.Z (CLOCK_slo___n64878), .A (n_6_4));
INV_X1 i_6_1_1663 (.ZN (n_6_2704), .A (n_6_1_879));
AOI222_X2 i_6_1_1662 (.ZN (n_6_1_878), .A1 (n_6_391), .A2 (n_6_1_904), .B1 (n_6_423)
    , .B2 (n_6_1_905), .C1 (n_6_2735), .C2 (CLOCK_sgo__n46934));
INV_X2 i_6_1_1661 (.ZN (n_6_2703), .A (n_6_1_878));
NAND2_X1 slo__sro_c13578 (.ZN (slo__sro_n12410), .A1 (n_6_2809), .A2 (n_6_1_973));
INV_X2 i_6_1_1659 (.ZN (n_6_2702), .A (n_6_1_877));
NAND2_X1 slo__sro_c13471 (.ZN (slo__sro_n12329), .A1 (n_6_2771), .A2 (CLOCK_sgo__n46937));
INV_X1 i_6_1_1657 (.ZN (n_6_2701), .A (slo__sro_n31816));
INV_X1 CLOCK_slo__sro_c56471 (.ZN (CLOCK_slo__sro_n51604), .A (slo__sro_n18951));
AOI21_X1 CLOCK_slo__sro_c54025 (.ZN (slo__sro_n9559), .A (CLOCK_slo__sro_n49402), .B1 (n_6_1320), .B2 (slo___n43257));
AOI222_X2 i_6_1_1654 (.ZN (CLOCK_sgo__n47094), .A1 (n_6_387), .A2 (n_6_1_904), .B1 (n_6_419)
    , .B2 (n_6_1_905), .C1 (n_6_2731), .C2 (CLOCK_sgo__n46934));
NAND2_X1 CLOCK_sgo__sro_c51476 (.ZN (CLOCK_sgo__sro_n47246), .A1 (slo___n13213), .A2 (n_6_1_168));
AOI222_X2 i_6_1_1652 (.ZN (n_6_1_873), .A1 (n_6_386), .A2 (n_6_1_904), .B1 (n_6_418)
    , .B2 (n_6_1_905), .C1 (n_6_2730), .C2 (CLOCK_sgo__n46934));
INV_X2 i_6_1_1651 (.ZN (n_6_2698), .A (n_6_1_873));
AND2_X1 slo__sro_c42822 (.ZN (slo__sro_n38699), .A1 (n_6_2382), .A2 (n_6_1_483));
INV_X1 CLOCK_slo__sro_c58030 (.ZN (CLOCK_slo__sro_n52917), .A (n_6_1_167));
INV_X1 CLOCK_slo__sro_c61541 (.ZN (CLOCK_slo__sro_n55890), .A (slo__sro_n11872));
INV_X2 i_6_1_1647 (.ZN (n_6_2696), .A (n_6_1_871));
NOR2_X4 i_6_1_1646 (.ZN (sgo__n594), .A1 (n_6_1_1123), .A2 (Multiplicand[7]));
NOR2_X4 i_6_1_1645 (.ZN (sgo__n607), .A1 (Multiplicand[8]), .A2 (n_6_1_1122));
NOR2_X4 i_6_1_1644 (.ZN (n_6_1_868), .A1 (n_6_1_870), .A2 (n_6_1_869));
AND2_X1 i_6_1_1643 (.ZN (n_6_1_867), .A1 (n_6_2726), .A2 (n_6_1_868));
AOI221_X2 i_6_1_1642 (.ZN (n_6_1_866), .A (n_6_1_867), .B1 (n_6_478), .B2 (n_6_1_869)
    , .C1 (n_6_510), .C2 (n_6_1_870));
INV_X1 i_6_1_1641 (.ZN (n_6_2695), .A (n_6_1_866));
AOI221_X1 i_6_1_1640 (.ZN (n_6_1_865), .A (n_6_1_867), .B1 (n_6_477), .B2 (n_6_1_869)
    , .C1 (n_6_509), .C2 (n_6_1_870));
INV_X1 i_6_1_1639 (.ZN (n_6_2694), .A (n_6_1_865));
NAND2_X1 slo__sro_c11416 (.ZN (slo__sro_n10561), .A1 (n_6_1818), .A2 (n_6_1_134));
INV_X1 i_6_1_1637 (.ZN (n_6_2693), .A (n_6_1_864));
NAND2_X1 slo__sro_c4464 (.ZN (slo__sro_n4288), .A1 (n_6_1_378), .A2 (n_6_2273));
INV_X1 i_6_1_1635 (.ZN (n_6_2692), .A (slo__sro_n4244));
AOI222_X2 i_6_1_1634 (.ZN (n_6_1_862), .A1 (n_6_506), .A2 (n_6_1_870), .B1 (n_6_474)
    , .B2 (n_6_1_869), .C1 (n_6_2723), .C2 (n_6_1_868));
INV_X1 CLOCK_sgo__sro_c52113 (.ZN (CLOCK_sgo__sro_n47762), .A (slo__sro_n20147));
AOI222_X2 i_6_1_1632 (.ZN (n_6_1_861), .A1 (n_6_505), .A2 (n_6_1_870), .B1 (n_6_473)
    , .B2 (n_6_1_869), .C1 (n_6_2722), .C2 (n_6_1_868));
INV_X1 i_6_1_1631 (.ZN (n_6_2690), .A (n_6_1_861));
BUF_X32 drc_ipo_c29979 (.Z (drc_ipo_n26602), .A (Multiplier[7]));
INV_X4 i_6_1_1629 (.ZN (n_6_2689), .A (CLOCK_slo__sro_n49602));
NAND2_X1 slo__sro_c8883 (.ZN (slo__sro_n8311), .A1 (n_6_2630), .A2 (n_6_1_763));
INV_X2 i_6_1_1627 (.ZN (n_6_2688), .A (slo__sro_n8294));
AOI222_X2 i_6_1_1626 (.ZN (slo__n26896), .A1 (n_6_502), .A2 (n_6_1_870), .B1 (n_6_470)
    , .B2 (n_6_1_869), .C1 (slo__n16557), .C2 (n_6_1_868));
INV_X1 slo__sro_c30282 (.ZN (slo__sro_n26911), .A (slo__sro_n26912));
AOI222_X2 i_6_1_1624 (.ZN (n_6_1_857), .A1 (n_6_501), .A2 (n_6_1_870), .B1 (n_6_469)
    , .B2 (n_6_1_869), .C1 (n_6_2718), .C2 (n_6_1_868));
INV_X2 i_6_1_1623 (.ZN (n_6_2686), .A (n_6_1_857));
NAND2_X1 slo__sro_c8199 (.ZN (slo__sro_n7692), .A1 (n_6_2463), .A2 (n_6_1_588));
INV_X4 i_6_1_1621 (.ZN (n_6_2685), .A (slo__sro_n20845));
NOR2_X1 slo__sro_c23025 (.ZN (slo__sro_n19998), .A1 (slo__sro_n20000), .A2 (slo__sro_n19999));
INV_X2 i_6_1_1619 (.ZN (n_6_2684), .A (slo__sro_n19894));
AND2_X1 slo__sro_c9169 (.ZN (slo__sro_n8559), .A1 (n_6_2567), .A2 (n_6_1_693));
INV_X1 i_6_1_1617 (.ZN (n_6_2683), .A (slo__sro_n8488));
AOI222_X2 slo__sro_c41003 (.ZN (n_6_1_1030), .A1 (n_6_179), .A2 (n_6_1_1045), .B1 (n_6_147)
    , .B2 (n_6_1_1044), .C1 (n_6_2871), .C2 (CLOCK_sgo__n46945));
INV_X2 i_6_1_1615 (.ZN (n_6_2682), .A (slo__sro_n37092));
NAND2_X2 CLOCK_slo__sro_c54228 (.ZN (CLOCK_slo__sro_n49604), .A1 (n_6_472), .A2 (n_6_1_869));
INV_X2 i_6_1_1613 (.ZN (n_6_2681), .A (CLOCK_slo__sro_n49426));
INV_X1 slo__sro_c33682 (.ZN (slo__sro_n30146), .A (CLOCK_sgo__n46934));
INV_X4 i_6_1_1611 (.ZN (n_6_2680), .A (n_6_1_851));
NAND2_X1 slo__sro_c41455 (.ZN (slo__sro_n37541), .A1 (n_6_518), .A2 (n_6_1_834));
INV_X1 i_6_1_1609 (.ZN (n_6_2679), .A (slo__sro_n37482));
AOI21_X1 slo__sro_c41087 (.ZN (slo__sro_n37221), .A (slo__sro_n37222), .B1 (n_6_124), .B2 (n_6_1_1080));
INV_X2 i_6_1_1607 (.ZN (n_6_2678), .A (n_6_1_849));
NAND2_X1 slo__sro_c40465 (.ZN (slo__sro_n36684), .A1 (n_6_2535), .A2 (n_6_1_658));
INV_X1 i_6_1_1605 (.ZN (n_6_2677), .A (CLOCK_slo__sro_n50400));
AOI221_X2 slo__sro_c37934 (.ZN (slo__sro_n34317), .A (slo__sro_n27159), .B1 (n_6_1914)
    , .B2 (n_6_1_100), .C1 (n_6_1882), .C2 (CLOCK_sgo__n48011));
INV_X2 i_6_1_1603 (.ZN (n_6_2676), .A (slo__sro_n33562));
NAND2_X1 CLOCK_slo__sro_c68588 (.ZN (CLOCK_slo__sro_n61784), .A1 (CLOCK_slo__sro_n61785), .A2 (CLOCK_slo__sro_n61786));
INV_X2 i_6_1_1601 (.ZN (n_6_2675), .A (slo__sro_n34126));
NAND2_X1 slo__sro_c9436 (.ZN (slo__sro_n8776), .A1 (slo__sro_n8777), .A2 (slo__sro_n8778));
NAND2_X1 CLOCK_slo__sro_c53531 (.ZN (CLOCK_slo__sro_n48977), .A1 (n_6_1803), .A2 (n_6_1_134));
INV_X2 slo__c16222 (.ZN (slo__n14603), .A (slo__sro_n8900));
INV_X1 i_6_1_1597 (.ZN (n_6_2673), .A (CLOCK_slo__sro_n59126));
AOI21_X1 slo__sro_c8441 (.ZN (slo__sro_n7910), .A (slo__sro_n7911), .B1 (n_6_628), .B2 (n_6_1_800));
INV_X2 i_6_1_1595 (.ZN (n_6_2672), .A (slo__sro_n7898));
NAND2_X1 slo__sro_c7250 (.ZN (slo__sro_n6829), .A1 (n_6_1260), .A2 (slo___n23274));
AOI21_X2 CLOCK_slo__sro_c71929 (.ZN (CLOCK_slo__sro_n64636), .A (CLOCK_slo__sro_n64637)
    , .B1 (n_6_1864), .B2 (CLOCK_sgo__n48011));
BUF_X32 drc_ipo_c29982 (.Z (drc_ipo_n26607), .A (Multiplier[12]));
INV_X2 i_6_1_1591 (.ZN (n_6_2670), .A (CLOCK_slo__sro_n48634));
NAND2_X1 slo__sro_c16917 (.ZN (slo__sro_n15200), .A1 (n_6_2650), .A2 (n_6_1_798));
NOR2_X1 CLOCK_slo__sro_c53218 (.ZN (CLOCK_slo__sro_n48698), .A1 (slo__sro_n9469), .A2 (CLOCK_slo__sro_n48699));
AOI21_X2 slo__sro_c12065 (.ZN (n_6_1_456), .A (slo__sro_n11124), .B1 (n_6_1189), .B2 (slo___n23466));
INV_X2 i_6_1_1587 (.ZN (n_6_2668), .A (n_6_1_839));
AND2_X1 slo__sro_c5006 (.ZN (slo__sro_n4775), .A1 (n_6_2409), .A2 (n_6_1_518));
INV_X4 i_6_1_1585 (.ZN (n_6_2667), .A (slo__sro_n4750));
NAND2_X1 CLOCK_slo__sro_c55281 (.ZN (CLOCK_slo__sro_n50547), .A1 (n_6_2433), .A2 (n_6_1_553));
INV_X1 i_6_1_1583 (.ZN (n_6_2666), .A (slo__sro_n6955));
AOI222_X1 i_6_1_1582 (.ZN (n_6_1_836), .A1 (n_6_448), .A2 (n_6_1_869), .B1 (n_6_480)
    , .B2 (n_6_1_870), .C1 (slo__n32451), .C2 (n_6_1_868));
INV_X1 i_6_1_1581 (.ZN (n_6_2665), .A (n_6_1_836));
NOR2_X4 i_6_1_1580 (.ZN (sgo__n566), .A1 (n_6_1_1124), .A2 (Multiplicand[8]));
NOR2_X4 i_6_1_1579 (.ZN (sgo__n577), .A1 (Multiplicand[9]), .A2 (n_6_1_1123));
NOR2_X4 i_6_1_1578 (.ZN (CLOCK_sgo__n46922), .A1 (n_6_1_835), .A2 (n_6_1_834));
AND2_X1 i_6_1_1577 (.ZN (n_6_1_832), .A1 (n_6_2695), .A2 (CLOCK_sgo__n46922));
AOI221_X1 i_6_1_1576 (.ZN (n_6_1_831), .A (n_6_1_832), .B1 (n_6_542), .B2 (n_6_1_834)
    , .C1 (n_6_574), .C2 (n_6_1_835));
INV_X1 i_6_1_1575 (.ZN (n_6_2664), .A (n_6_1_831));
AOI221_X2 i_6_1_1574 (.ZN (n_6_1_830), .A (n_6_1_832), .B1 (n_6_541), .B2 (n_6_1_834)
    , .C1 (n_6_573), .C2 (n_6_1_835));
INV_X2 i_6_1_1573 (.ZN (n_6_2663), .A (n_6_1_830));
NAND2_X1 slo__sro_c13777 (.ZN (slo__sro_n12571), .A1 (n_6_1_413), .A2 (n_6_2318));
INV_X2 i_6_1_1571 (.ZN (n_6_2662), .A (n_6_1_829));
AOI222_X2 i_6_1_1570 (.ZN (n_6_1_828), .A1 (n_6_571), .A2 (n_6_1_835), .B1 (n_6_539)
    , .B2 (n_6_1_834), .C1 (n_6_2693), .C2 (CLOCK_sgo__n46922));
INV_X1 i_6_1_1569 (.ZN (n_6_2661), .A (n_6_1_828));
AOI21_X1 CLOCK_slo__sro_c62452 (.ZN (CLOCK_slo__sro_n56609), .A (slo__sro_n20923)
    , .B1 (n_6_182), .B2 (n_6_1_1045));
INV_X1 i_6_1_1567 (.ZN (n_6_2660), .A (n_6_1_827));
AOI222_X2 slo__sro_c12341 (.ZN (n_6_1_714), .A1 (n_6_722), .A2 (n_6_1_729), .B1 (n_6_754)
    , .B2 (n_6_1_730), .C1 (n_6_2591), .C2 (n_6_1_728));
INV_X1 i_6_1_1565 (.ZN (n_6_2659), .A (slo__sro_n11215));
AOI222_X2 slo__sro_c8076 (.ZN (slo__sro_n7583), .A1 (n_6_438), .A2 (n_6_1_905), .B1 (n_6_406)
    , .B2 (n_6_1_904), .C1 (n_6_2750), .C2 (CLOCK_sgo__n46934));
INV_X1 i_6_1_1563 (.ZN (n_6_2658), .A (n_6_1_825));
NAND2_X1 CLOCK_sgo__sro_c51910 (.ZN (CLOCK_sgo__sro_n47604), .A1 (n_6_1_133), .A2 (n_6_2068));
INV_X1 i_6_1_1561 (.ZN (n_6_2657), .A (n_6_1_824));
AOI21_X1 CLOCK_slo__sro_c67394 (.ZN (CLOCK_slo__sro_n60680), .A (slo__sro_n8978), .B1 (n_6_346), .B2 (n_6_1_939));
INV_X2 i_6_1_1559 (.ZN (n_6_2656), .A (CLOCK_slo__sro_n56376));
NAND2_X1 slo__sro_c9220 (.ZN (slo__sro_n8605), .A1 (slo__n13799), .A2 (n_6_2885));
INV_X1 i_6_1_1557 (.ZN (slo___n19273), .A (slo__sro_n30031));
AND2_X1 CLOCK_slo__sro_c64864 (.ZN (CLOCK_slo__sro_n58451), .A1 (n_6_2884), .A2 (slo__n13799));
INV_X2 i_6_1_1555 (.ZN (slo___n19182), .A (slo__sro_n8500));
AOI222_X2 i_6_1_1554 (.ZN (n_6_1_820), .A1 (n_6_563), .A2 (n_6_1_835), .B1 (n_6_531)
    , .B2 (n_6_1_834), .C1 (n_6_2685), .C2 (CLOCK_sgo__n46922));
INV_X2 i_6_1_1553 (.ZN (n_6_2653), .A (n_6_1_820));
AOI21_X1 slo__sro_c9437 (.ZN (n_6_1_1021), .A (slo__sro_n8776), .B1 (n_6_138), .B2 (n_6_1_1044));
INV_X1 i_6_1_1551 (.ZN (n_6_2652), .A (n_6_1_819));
INV_X1 slo__sro_c22996 (.ZN (slo__sro_n19973), .A (n_6_2461));
INV_X2 i_6_1_1549 (.ZN (n_6_2651), .A (slo__sro_n19805));
NAND2_X1 slo__sro_c12448 (.ZN (slo__sro_n11438), .A1 (n_6_2393), .A2 (n_6_1_518));
INV_X1 i_6_1_1547 (.ZN (n_6_2650), .A (CLOCK_slo__sro_n60275));
NAND2_X1 slo__sro_c5551 (.ZN (slo__sro_n5285), .A1 (n_6_2678), .A2 (CLOCK_sgo__n46922));
INV_X1 i_6_1_1545 (.ZN (n_6_2649), .A (CLOCK_slo__sro_n51643));
AND2_X1 CLOCK_slo__sro_c62633 (.ZN (CLOCK_slo__sro_n56757), .A1 (n_6_562), .A2 (n_6_1_835));
INV_X2 i_6_1_1543 (.ZN (n_6_2648), .A (n_6_1_815));
NAND2_X1 slo__sro_c46315 (.ZN (slo__sro_n41809), .A1 (n_6_1753), .A2 (n_6_1_169));
INV_X2 i_6_1_1541 (.ZN (n_6_2647), .A (slo__sro_n7219));
BUF_X1 slo__c5578 (.Z (spw__n66887), .A (sgo__n1271));
INV_X2 i_6_1_1539 (.ZN (n_6_2646), .A (n_6_1_813));
AOI21_X1 CLOCK_slo__sro_c58227 (.ZN (n_6_1_1055), .A (CLOCK_slo__sro_n53078), .B1 (n_6_73), .B2 (n_6_1_1079));
INV_X1 i_6_1_1537 (.ZN (n_6_2645), .A (CLOCK_slo__sro_n53015));
AOI222_X1 i_6_1_1536 (.ZN (n_6_1_811), .A1 (n_6_522), .A2 (n_6_1_834), .B1 (n_6_554)
    , .B2 (n_6_1_835), .C1 (n_6_2676), .C2 (CLOCK_sgo__n46922));
INV_X1 i_6_1_1535 (.ZN (n_6_2644), .A (n_6_1_811));
NAND2_X1 slo__sro_c6611 (.ZN (slo__sro_n6242), .A1 (n_6_2703), .A2 (n_6_1_868));
INV_X1 i_6_1_1533 (.ZN (slo___n15116), .A (slo__sro_n6229));
AOI222_X1 CLOCK_slo__sro_c63179 (.ZN (n_6_1_919), .A1 (n_6_365), .A2 (n_6_1_940), .B1 (n_6_333)
    , .B2 (n_6_1_939), .C1 (n_6_2772), .C2 (CLOCK_sgo__n46937));
INV_X2 i_6_1_1531 (.ZN (n_6_2642), .A (n_6_1_809));
AOI222_X2 i_6_1_1530 (.ZN (n_6_1_808), .A1 (n_6_519), .A2 (n_6_1_834), .B1 (n_6_551)
    , .B2 (n_6_1_835), .C1 (n_6_2673), .C2 (CLOCK_sgo__n46922));
INV_X2 i_6_1_1529 (.ZN (n_6_2641), .A (n_6_1_808));
NAND2_X1 slo__sro_c33379 (.ZN (slo__sro_n29860), .A1 (slo__n30795), .A2 (n_6_1_203));
INV_X4 i_6_1_1527 (.ZN (n_6_2640), .A (slo__sro_n37539));
AND2_X2 CLOCK_slo__sro_c61696 (.ZN (CLOCK_slo__sro_n56009), .A1 (n_6_89), .A2 (n_6_1_1079));
INV_X2 i_6_1_1525 (.ZN (n_6_2639), .A (n_6_1_806));
NAND2_X1 slo__sro_c21156 (.ZN (slo__sro_n18492), .A1 (n_6_2702), .A2 (n_6_1_868));
INV_X1 i_6_1_1523 (.ZN (n_6_2638), .A (CLOCK_slo__sro_n56126));
NAND2_X1 slo__sro_c38397 (.ZN (slo__sro_n34758), .A1 (n_6_2208), .A2 (n_6_1_308));
INV_X2 i_6_1_1521 (.ZN (n_6_2637), .A (slo__sro_n15043));
AOI222_X2 i_6_1_1520 (.ZN (n_6_1_803), .A1 (n_6_514), .A2 (n_6_1_834), .B1 (n_6_546)
    , .B2 (n_6_1_835), .C1 (n_6_2668), .C2 (CLOCK_sgo__n46922));
INV_X2 i_6_1_1519 (.ZN (n_6_2636), .A (n_6_1_803));
INV_X1 CLOCK_slo__sro_c62808 (.ZN (CLOCK_slo__sro_n56896), .A (slo__sro_n15796));
INV_X1 i_6_1_1517 (.ZN (n_6_2635), .A (n_6_1_802));
AOI222_X1 i_6_1_1516 (.ZN (spt__n66327), .A1 (n_6_512), .A2 (n_6_1_834), .B1 (n_6_544)
    , .B2 (n_6_1_835), .C1 (n_6_2666), .C2 (CLOCK_sgo__n46922));
INV_X2 i_6_1_1515 (.ZN (n_6_2634), .A (n_6_1_801));
NOR2_X4 i_6_1_1514 (.ZN (sgo__n544), .A1 (n_6_1_1125), .A2 (Multiplicand[9]));
NOR2_X4 i_6_1_1513 (.ZN (sgo__n553), .A1 (Multiplicand[10]), .A2 (n_6_1_1124));
NOR2_X4 i_6_1_1512 (.ZN (n_6_1_798), .A1 (n_6_1_800), .A2 (n_6_1_799));
AND2_X1 i_6_1_1511 (.ZN (n_6_1_797), .A1 (n_6_2664), .A2 (n_6_1_798));
AOI221_X1 i_6_1_1510 (.ZN (n_6_1_796), .A (n_6_1_797), .B1 (n_6_606), .B2 (n_6_1_799)
    , .C1 (n_6_638), .C2 (n_6_1_800));
INV_X1 i_6_1_1509 (.ZN (n_6_2633), .A (n_6_1_796));
AOI221_X1 i_6_1_1508 (.ZN (n_6_1_795), .A (n_6_1_797), .B1 (n_6_605), .B2 (n_6_1_799)
    , .C1 (n_6_637), .C2 (n_6_1_800));
INV_X1 i_6_1_1507 (.ZN (n_6_2632), .A (n_6_1_795));
NAND2_X1 slo__sro_c13762 (.ZN (slo__sro_n12557), .A1 (n_6_540), .A2 (n_6_1_834));
INV_X2 i_6_1_1505 (.ZN (n_6_2631), .A (n_6_1_794));
AND2_X1 slo__sro_c11366 (.ZN (slo__sro_n10518), .A1 (n_6_2725), .A2 (n_6_1_868));
INV_X2 i_6_1_1503 (.ZN (n_6_2630), .A (n_6_1_793));
AOI222_X2 i_6_1_1502 (.ZN (n_6_1_792), .A1 (n_6_634), .A2 (n_6_1_800), .B1 (n_6_602)
    , .B2 (n_6_1_799), .C1 (n_6_2661), .C2 (n_6_1_798));
INV_X1 i_6_1_1501 (.ZN (n_6_2629), .A (n_6_1_792));
NAND2_X1 slo__sro_c4403 (.ZN (slo__sro_n4233), .A1 (n_6_2563), .A2 (n_6_1_693));
INV_X1 i_6_1_1499 (.ZN (n_6_2628), .A (n_6_1_791));
INV_X1 CLOCK_slo__sro_c58324 (.ZN (CLOCK_slo__sro_n53159), .A (slo__sro_n30922));
INV_X2 i_6_1_1497 (.ZN (n_6_2627), .A (n_6_1_790));
AOI222_X2 i_6_1_1496 (.ZN (n_6_1_789), .A1 (n_6_631), .A2 (n_6_1_800), .B1 (n_6_599)
    , .B2 (n_6_1_799), .C1 (n_6_2658), .C2 (n_6_1_798));
INV_X1 i_6_1_1495 (.ZN (n_6_2626), .A (n_6_1_789));
AOI21_X2 slo__sro_c8870 (.ZN (slo__sro_n8294), .A (slo__sro_n8295), .B1 (n_6_503), .B2 (n_6_1_870));
INV_X2 i_6_1_1493 (.ZN (n_6_2625), .A (n_6_1_788));
INV_X2 opt_ipo_c29621 (.ZN (opt_ipo_n26244), .A (slo__sro_n13700));
INV_X1 i_6_1_1491 (.ZN (slo___n12846), .A (slo__sro_n21940));
NAND2_X1 slo__sro_c8472 (.ZN (slo__sro_n7947), .A1 (n_6_2907), .A2 (slo__n13799));
INV_X2 i_6_1_1489 (.ZN (n_6_2623), .A (slo__sro_n7910));
INV_X1 slo__c22195 (.ZN (slo__n19260), .A (slo__sro_n7944));
INV_X1 i_6_1_1487 (.ZN (n_6_2622), .A (slo__sro_n19076));
AND2_X1 slo__sro_c7049 (.ZN (slo__sro_n6654), .A1 (n_6_2300), .A2 (n_6_1_413));
INV_X2 i_6_1_1485 (.ZN (n_6_2621), .A (slo__sro_n20817));
INV_X1 slo___L2_c4_c14397 (.ZN (n_6_2070), .A (slo___n13099));
NAND2_X1 slo__sro_c33403 (.ZN (slo__sro_n29881), .A1 (n_6_482), .A2 (n_6_1_870));
NAND2_X1 slo__sro_c12064 (.ZN (slo__sro_n11124), .A1 (slo__sro_n11125), .A2 (slo__sro_n11126));
NAND2_X1 CLOCK_slo__sro_c55754 (.ZN (CLOCK_slo__sro_n50976), .A1 (n_6_2618), .A2 (n_6_1_763));
AOI222_X1 slo__sro_c17125 (.ZN (n_6_1_875), .A1 (n_6_420), .A2 (n_6_1_905), .B1 (n_6_388)
    , .B2 (n_6_1_904), .C1 (n_6_2732), .C2 (CLOCK_sgo__n46934));
INV_X2 i_6_1_1479 (.ZN (n_6_2618), .A (CLOCK_slo__sro_n51723));
NAND2_X1 CLOCK_slo__sro_c53834 (.ZN (CLOCK_slo__sro_n49244), .A1 (n_6_2412), .A2 (n_6_1_518));
INV_X2 i_6_1_1477 (.ZN (n_6_2617), .A (CLOCK_slo__sro_n49188));
INV_X4 slo__c15598 (.ZN (slo__n14062), .A (n_6_1_699));
INV_X1 i_6_1_1475 (.ZN (n_6_2616), .A (n_6_1_779));
NAND2_X1 slo__sro_c18206 (.ZN (slo__sro_n16217), .A1 (n_6_168), .A2 (n_6_1_1045));
INV_X1 i_6_1_1473 (.ZN (n_6_2615), .A (slo__sro_n16180));
AOI222_X2 i_6_1_1472 (.ZN (n_6_1_777), .A1 (n_6_587), .A2 (n_6_1_799), .B1 (n_6_619)
    , .B2 (n_6_1_800), .C1 (n_6_2646), .C2 (n_6_1_798));
INV_X2 i_6_1_1471 (.ZN (n_6_2614), .A (n_6_1_777));
INV_X1 slo__sro_c11190 (.ZN (slo__sro_n10380), .A (n_6_2755));
INV_X1 i_6_1_1469 (.ZN (n_6_2613), .A (slo__sro_n10270));
BUF_X16 drc_ipo_c29967 (.Z (drc_ipo_n26590), .A (n_6_9));
INV_X2 i_6_1_1467 (.ZN (n_6_2612), .A (n_6_1_775));
NAND2_X1 CLOCK_slo__sro_c69381 (.ZN (CLOCK_slo__sro_n62489), .A1 (n_6_458), .A2 (n_6_1_869));
INV_X2 i_6_1_1465 (.ZN (n_6_2611), .A (slo__sro_n32026));
NAND2_X1 slo__sro_c25142 (.ZN (slo__sro_n21942), .A1 (n_6_629), .A2 (n_6_1_800));
INV_X2 i_6_1_1463 (.ZN (n_6_2610), .A (n_6_1_773));
AOI221_X2 slo__sro_c6000 (.ZN (slo__sro_n5678), .A (slo__sro_n5679), .B1 (n_6_1166)
    , .B2 (slo___n23364), .C1 (n_6_1198), .C2 (slo___n23466));
INV_X1 i_6_1_1461 (.ZN (n_6_2609), .A (slo__sro_n5416));
NAND2_X1 slo__sro_c35469 (.ZN (slo__sro_n31832), .A1 (n_6_2831), .A2 (CLOCK_sgo__n46950));
INV_X4 i_6_1_1459 (.ZN (n_6_2608), .A (slo__sro_n12110));
NAND2_X1 slo__sro_c31974 (.ZN (slo__sro_n28526), .A1 (n_6_2585), .A2 (n_6_1_728));
INV_X2 i_6_1_1457 (.ZN (n_6_2607), .A (n_6_1_770));
INV_X1 CLOCK_slo__sro_c65144 (.ZN (CLOCK_slo__sro_n58700), .A (slo__sro_n40960));
NAND2_X1 CLOCK_slo__sro_c64711 (.ZN (CLOCK_slo__sro_n58341), .A1 (CLOCK_slo__sro_n58342), .A2 (CLOCK_slo__sro_n58343));
AOI21_X2 slo__sro_c45536 (.ZN (slo__sro_n41060), .A (slo__sro_n19450), .B1 (n_6_791), .B2 (n_6_1_694));
INV_X2 i_6_1_1453 (.ZN (CLOCK_slo___n54911), .A (slo__sro_n40959));
INV_X1 CLOCK_slo__c61039 (.ZN (CLOCK_slo__n55465), .A (n_6_1_347));
INV_X2 i_6_1_1451 (.ZN (n_6_2604), .A (n_6_1_767));
AOI222_X1 i_6_1_1450 (.ZN (n_6_1_766), .A1 (n_6_576), .A2 (n_6_1_799), .B1 (n_6_608)
    , .B2 (n_6_1_800), .C1 (n_6_2635), .C2 (n_6_1_798));
INV_X1 i_6_1_1449 (.ZN (CLOCK_slo___n64354), .A (n_6_1_766));
NOR2_X1 i_6_1_1448 (.ZN (sgo__n521), .A1 (n_6_1_1126), .A2 (Multiplicand[10]));
NOR2_X4 i_6_1_1447 (.ZN (sgo__n535), .A1 (Multiplicand[11]), .A2 (n_6_1_1125));
NOR2_X4 i_6_1_1446 (.ZN (n_6_1_763), .A1 (n_6_1_765), .A2 (n_6_1_764));
AND2_X1 i_6_1_1445 (.ZN (n_6_1_762), .A1 (n_6_2633), .A2 (n_6_1_763));
AOI221_X2 i_6_1_1444 (.ZN (n_6_1_761), .A (n_6_1_762), .B1 (n_6_670), .B2 (n_6_1_764)
    , .C1 (n_6_702), .C2 (n_6_1_765));
INV_X2 i_6_1_1443 (.ZN (n_6_2602), .A (n_6_1_761));
AOI221_X2 i_6_1_1442 (.ZN (n_6_1_760), .A (n_6_1_762), .B1 (n_6_669), .B2 (n_6_1_764)
    , .C1 (n_6_701), .C2 (n_6_1_765));
INV_X1 i_6_1_1441 (.ZN (n_6_2601), .A (n_6_1_760));
NAND2_X1 slo__sro_c13221 (.ZN (slo__sro_n12112), .A1 (n_6_613), .A2 (n_6_1_800));
INV_X2 i_6_1_1439 (.ZN (n_6_2600), .A (n_6_1_759));
NAND2_X1 slo__sro_c10729 (.ZN (slo__sro_n9979), .A1 (n_6_2442), .A2 (n_6_1_553));
INV_X2 slo__c40090 (.ZN (slo__n36350), .A (slo__sro_n12647));
BUF_X32 drc_ipo_c29966 (.Z (drc_ipo_n26589), .A (n_6_11));
NAND2_X1 slo__sro_c33191 (.ZN (slo__sro_n29676), .A1 (n_6_270), .A2 (n_6_1_974));
AOI222_X2 slo__sro_c41147 (.ZN (n_6_1_635), .A1 (n_6_841), .A2 (slo___n23463), .B1 (n_6_873)
    , .B2 (n_6_1_660), .C1 (n_6_2520), .C2 (n_6_1_658));
INV_X1 i_6_1_1433 (.ZN (n_6_2597), .A (n_6_1_756));
AOI222_X2 i_6_1_1432 (.ZN (n_6_1_755), .A1 (n_6_696), .A2 (n_6_1_765), .B1 (n_6_664)
    , .B2 (n_6_1_764), .C1 (n_6_2628), .C2 (n_6_1_763));
INV_X2 i_6_1_1431 (.ZN (n_6_2596), .A (n_6_1_755));
INV_X2 i_6_1_1429 (.ZN (n_6_2595), .A (n_6_1_754));
AOI21_X4 slo__sro_c25342 (.ZN (slo__sro_n22134), .A (slo__sro_n13318), .B1 (n_6_1623), .B2 (slo___n23215));
INV_X4 i_6_1_1427 (.ZN (n_6_2594), .A (slo__sro_n22110));
NAND2_X1 slo__sro_c38853 (.ZN (slo__sro_n35199), .A1 (n_6_2827), .A2 (CLOCK_sgo__n46950));
INV_X1 i_6_1_1425 (.ZN (n_6_2593), .A (slo__sro_n35183));
NAND2_X1 slo__sro_c32551 (.ZN (slo__sro_n29069), .A1 (n_6_2050), .A2 (n_6_1_133));
INV_X4 i_6_1_1423 (.ZN (n_6_2592), .A (slo__sro_n28774));
INV_X1 CLOCK_slo__c61574 (.ZN (CLOCK_slo__n55908), .A (slo__sro_n4244));
INV_X2 i_6_1_1421 (.ZN (n_6_2591), .A (CLOCK_slo__sro_n55784));
NAND2_X1 CLOCK_slo__sro_c68487 (.ZN (CLOCK_slo__sro_n61696), .A1 (CLOCK_slo__sro_n61697), .A2 (CLOCK_slo__sro_n61698));
INV_X2 i_6_1_1419 (.ZN (n_6_2590), .A (n_6_1_749));
AOI222_X2 i_6_1_1418 (.ZN (n_6_1_748), .A1 (n_6_689), .A2 (n_6_1_765), .B1 (n_6_657)
    , .B2 (n_6_1_764), .C1 (n_6_2621), .C2 (n_6_1_763));
INV_X2 i_6_1_1417 (.ZN (n_6_2589), .A (n_6_1_748));
AND2_X1 CLOCK_slo__sro_c55932 (.ZN (CLOCK_slo__sro_n51133), .A1 (slo___n17886), .A2 (n_6_1_588));
INV_X2 i_6_1_1415 (.ZN (n_6_2588), .A (CLOCK_slo__sro_n51092));
NAND2_X1 slo__sro_c11067 (.ZN (slo__sro_n10272), .A1 (n_6_618), .A2 (n_6_1_800));
INV_X2 i_6_1_1413 (.ZN (n_6_2587), .A (slo__sro_n34034));
NAND2_X1 CLOCK_slo__sro_c55773 (.ZN (CLOCK_slo__sro_n50987), .A1 (n_6_1532), .A2 (slo___n23247));
INV_X2 i_6_1_1411 (.ZN (n_6_2586), .A (n_6_1_745));
NAND2_X1 slo__sro_c31104 (.ZN (slo__sro_n27690), .A1 (slo__sro_n27691), .A2 (slo__sro_n10080));
INV_X2 i_6_1_1409 (.ZN (n_6_2585), .A (n_6_1_744));
AOI222_X2 i_6_1_1408 (.ZN (n_6_1_743), .A1 (n_6_652), .A2 (n_6_1_764), .B1 (n_6_684)
    , .B2 (n_6_1_765), .C1 (n_6_2616), .C2 (n_6_1_763));
INV_X2 i_6_1_1407 (.ZN (n_6_2584), .A (n_6_1_743));
BUF_X32 drc_ipo_c29980 (.Z (drc_ipo_n26605), .A (Multiplier[10]));
INV_X1 i_6_1_1405 (.ZN (n_6_2583), .A (CLOCK_slo__sro_n62823));
AND2_X1 slo__sro_c6340 (.ZN (slo__sro_n5988), .A1 (n_6_2487), .A2 (n_6_1_623));
INV_X2 i_6_1_1403 (.ZN (n_6_2582), .A (n_6_1_741));
AND2_X1 slo__sro_c8606 (.ZN (slo__sro_n8057), .A1 (n_6_1_757), .A2 (n_6_1_728));
INV_X1 i_6_1_1401 (.ZN (n_6_2581), .A (slo__sro_n27860));
BUF_X32 drc_ipo_c29961 (.Z (drc_ipo_n26584), .A (n_6_15));
AOI221_X2 CLOCK_slo__sro_c53320 (.ZN (CLOCK_slo__sro_n48784), .A (CLOCK_slo__sro_n48785)
    , .B1 (n_6_1498), .B2 (n_6_1_309), .C1 (n_6_1530), .C2 (slo___n23247));
NAND2_X1 slo__sro_c8440 (.ZN (slo__sro_n7911), .A1 (slo__sro_n7912), .A2 (slo__sro_n7913));
INV_X1 i_6_1_1397 (.ZN (slo___n13777), .A (slo__sro_n19436));
NAND2_X1 slo__sro_c16535 (.ZN (slo__sro_n14857), .A1 (n_6_2586), .A2 (n_6_1_728));
NAND2_X2 CLOCK_slo__sro_c54053 (.ZN (CLOCK_slo__sro_n49427), .A1 (CLOCK_slo__sro_n49428), .A2 (CLOCK_slo__sro_n49429));
NAND2_X1 slo__sro_c38839 (.ZN (slo__sro_n35186), .A1 (n_6_2625), .A2 (n_6_1_763));
INV_X1 i_6_1_1393 (.ZN (n_6_2577), .A (slo__sro_n35163));
INV_X1 slo__sro_c12490 (.ZN (slo__sro_n11473), .A (slo__sro_n11474));
INV_X2 i_6_1_1391 (.ZN (n_6_2576), .A (slo__sro_n37387));
NAND2_X1 slo__sro_c13220 (.ZN (slo__sro_n12113), .A1 (n_6_1_798), .A2 (n_6_2640));
NAND2_X2 CLOCK_slo__sro_c53836 (.ZN (CLOCK_slo__sro_n49242), .A1 (CLOCK_slo__sro_n49243), .A2 (CLOCK_slo__sro_n49244));
AOI222_X2 i_6_1_1388 (.ZN (n_6_1_733), .A1 (n_6_642), .A2 (n_6_1_764), .B1 (n_6_674)
    , .B2 (n_6_1_765), .C1 (opt_ipo_n44394), .C2 (n_6_1_763));
INV_X2 i_6_1_1387 (.ZN (n_6_2574), .A (n_6_1_733));
AOI222_X1 i_6_1_1386 (.ZN (n_6_1_732), .A1 (n_6_641), .A2 (n_6_1_764), .B1 (n_6_673)
    , .B2 (n_6_1_765), .C1 (CLOCK_slo___n54911), .C2 (n_6_1_763));
INV_X1 i_6_1_1385 (.ZN (n_6_2573), .A (n_6_1_732));
AOI222_X1 i_6_1_1384 (.ZN (n_6_1_731), .A1 (n_6_640), .A2 (n_6_1_764), .B1 (n_6_672)
    , .B2 (n_6_1_765), .C1 (n_6_2604), .C2 (n_6_1_763));
INV_X1 i_6_1_1383 (.ZN (spw__n67889), .A (n_6_1_731));
NOR2_X4 i_6_1_1382 (.ZN (sgo__n495), .A1 (n_6_1_1127), .A2 (Multiplicand[11]));
NOR2_X4 i_6_1_1381 (.ZN (sgo__n508), .A1 (Multiplicand[12]), .A2 (n_6_1_1126));
NOR2_X4 i_6_1_1380 (.ZN (n_6_1_728), .A1 (n_6_1_730), .A2 (n_6_1_729));
AND2_X1 i_6_1_1379 (.ZN (n_6_1_727), .A1 (n_6_2602), .A2 (n_6_1_728));
AOI221_X1 i_6_1_1378 (.ZN (n_6_1_726), .A (n_6_1_727), .B1 (n_6_734), .B2 (n_6_1_729)
    , .C1 (n_6_766), .C2 (n_6_1_730));
INV_X1 i_6_1_1377 (.ZN (n_6_2571), .A (n_6_1_726));
AOI221_X2 i_6_1_1376 (.ZN (n_6_1_725), .A (n_6_1_727), .B1 (n_6_733), .B2 (n_6_1_729)
    , .C1 (n_6_765), .C2 (n_6_1_730));
INV_X1 i_6_1_1375 (.ZN (n_6_2570), .A (n_6_1_725));
AOI222_X2 i_6_1_1374 (.ZN (n_6_1_724), .A1 (n_6_764), .A2 (n_6_1_730), .B1 (n_6_732)
    , .B2 (n_6_1_729), .C1 (n_6_2601), .C2 (n_6_1_728));
INV_X2 i_6_1_1373 (.ZN (n_6_2569), .A (n_6_1_724));
NAND2_X1 slo__sro_c9582 (.ZN (slo__sro_n8919), .A1 (n_6_1_693), .A2 (n_6_2545));
INV_X2 i_6_1_1371 (.ZN (n_6_2568), .A (n_6_1_723));
INV_X1 slo__sro_c10869 (.ZN (slo__sro_n10100), .A (n_6_2754));
INV_X1 i_6_1_1369 (.ZN (n_6_2567), .A (slo__sro_n27689));
NAND2_X1 slo__sro_c35859 (.ZN (slo__sro_n32203), .A1 (n_6_1754), .A2 (n_6_1_169));
INV_X4 i_6_1_1367 (.ZN (n_6_2566), .A (slo__sro_n27581));
NAND2_X1 slo__sro_c8592 (.ZN (slo__sro_n8047), .A1 (n_6_2617), .A2 (n_6_1_763));
INV_X2 i_6_1_1365 (.ZN (n_6_2565), .A (n_6_1_720));
INV_X1 slo__sro_c30904 (.ZN (slo__sro_n27500), .A (slo__sro_n27501));
INV_X1 i_6_1_1363 (.ZN (n_6_2564), .A (n_6_1_719));
NAND2_X1 slo__sro_c10849 (.ZN (slo__sro_n10080), .A1 (slo__n35732), .A2 (n_6_1_728));
INV_X2 i_6_1_1361 (.ZN (n_6_2563), .A (n_6_1_718));
AOI222_X2 i_6_1_1360 (.ZN (n_6_1_717), .A1 (n_6_757), .A2 (n_6_1_730), .B1 (n_6_725)
    , .B2 (n_6_1_729), .C1 (n_6_2594), .C2 (n_6_1_728));
INV_X1 i_6_1_1359 (.ZN (n_6_2562), .A (n_6_1_717));
AOI221_X1 slo__sro_c37469 (.ZN (slo__sro_n33788), .A (slo__sro_n33789), .B1 (n_6_810)
    , .B2 (n_6_1_695), .C1 (n_6_778), .C2 (n_6_1_694));
INV_X2 i_6_1_1357 (.ZN (n_6_2561), .A (slo__sro_n33706));
NAND2_X1 slo__sro_c13687 (.ZN (slo__sro_n12493), .A1 (n_6_2506), .A2 (n_6_1_623));
INV_X1 i_6_1_1355 (.ZN (n_6_2560), .A (slo__sro_n12465));
NAND2_X1 slo__sro_c12449 (.ZN (slo__sro_n11437), .A1 (n_6_1126), .A2 (slo___n23268));
INV_X2 i_6_1_1353 (.ZN (n_6_2559), .A (n_6_1_714));
NAND2_X1 slo__sro_c14191 (.ZN (slo__sro_n12926), .A1 (n_6_1_273), .A2 (n_6_2184));
INV_X2 i_6_1_1351 (.ZN (n_6_2558), .A (n_6_1_713));
AND2_X1 slo__sro_c16205 (.ZN (slo__sro_n14590), .A1 (n_6_2526), .A2 (n_6_1_658));
INV_X1 i_6_1_1349 (.ZN (n_6_2557), .A (n_6_1_712));
NAND2_X1 slo__sro_c22362 (.ZN (slo__sro_n19385), .A1 (n_6_1_973), .A2 (n_6_2816));
INV_X1 i_6_1_1347 (.ZN (n_6_2556), .A (n_6_1_711));
AOI221_X1 slo__sro_c8740 (.ZN (slo__n29395), .A (slo__sro_n8180), .B1 (n_6_986), .B2 (slo___n23232)
    , .C1 (n_6_1018), .C2 (slo___n23218));
INV_X4 i_6_1_1345 (.ZN (n_6_2555), .A (slo__sro_n7705));
AND2_X1 slo__sro_c16601 (.ZN (slo__sro_n14915), .A1 (n_6_2615), .A2 (n_6_1_763));
INV_X4 i_6_1_1343 (.ZN (n_6_2554), .A (slo__sro_n14854));
AOI222_X1 CLOCK_slo__sro_c58985 (.ZN (n_6_1_398), .A1 (n_6_1297), .A2 (n_6_1_414)
    , .B1 (n_6_1329), .B2 (slo___n43257), .C1 (n_6_2311), .C2 (n_6_1_413));
INV_X1 i_6_1_1341 (.ZN (n_6_2553), .A (slo__sro_n28523));
NAND2_X1 slo__sro_c5631 (.ZN (slo__sro_n5354), .A1 (n_6_2774), .A2 (CLOCK_sgo__n46937));
INV_X4 i_6_1_1339 (.ZN (n_6_2552), .A (n_6_1_707));
AOI222_X2 i_6_1_1338 (.ZN (n_6_1_706), .A1 (n_6_714), .A2 (n_6_1_729), .B1 (n_6_746)
    , .B2 (n_6_1_730), .C1 (n_6_2583), .C2 (n_6_1_728));
INV_X1 i_6_1_1337 (.ZN (n_6_2551), .A (n_6_1_706));
AOI21_X2 slo__sro_c16538 (.ZN (slo__sro_n14854), .A (slo__sro_n14855), .B1 (n_6_749), .B2 (n_6_1_730));
INV_X1 i_6_1_1335 (.ZN (slo___n17474), .A (CLOCK_slo__sro_n54647));
AOI222_X2 i_6_1_1334 (.ZN (n_6_1_704), .A1 (n_6_712), .A2 (n_6_1_729), .B1 (n_6_744)
    , .B2 (n_6_1_730), .C1 (n_6_2581), .C2 (n_6_1_728));
INV_X2 i_6_1_1333 (.ZN (n_6_2549), .A (n_6_1_704));
AOI222_X2 i_6_1_1332 (.ZN (n_6_1_703), .A1 (n_6_711), .A2 (n_6_1_729), .B1 (n_6_743)
    , .B2 (n_6_1_730), .C1 (CLOCK_opt_ipo_n46029), .C2 (n_6_1_728));
INV_X2 i_6_1_1331 (.ZN (n_6_2548), .A (n_6_1_703));
INV_X1 i_6_1_1329 (.ZN (n_6_2547), .A (slo__sro_n42331));
INV_X1 slo__sro_c13579 (.ZN (slo__sro_n12409), .A (slo__sro_n12410));
INV_X2 i_6_1_1327 (.ZN (n_6_2546), .A (slo__sro_n12255));
AOI222_X2 i_6_1_1326 (.ZN (n_6_1_700), .A1 (n_6_708), .A2 (n_6_1_729), .B1 (n_6_740)
    , .B2 (n_6_1_730), .C1 (n_6_2577), .C2 (n_6_1_728));
INV_X2 i_6_1_1325 (.ZN (n_6_2545), .A (n_6_1_700));
AOI221_X2 slo__sro_c38193 (.ZN (slo__sro_n34553), .A (slo__sro_n34554), .B1 (n_6_1561)
    , .B2 (n_6_1_274), .C1 (n_6_1593), .C2 (slo___n23244));
INV_X1 i_6_1_1323 (.ZN (n_6_2544), .A (n_6_1_699));
NAND2_X1 slo__sro_c25023 (.ZN (slo__sro_n21836), .A1 (n_6_2807), .A2 (n_6_1_973));
INV_X2 i_6_1_1321 (.ZN (n_6_2543), .A (slo__sro_n21676));
AOI222_X2 i_6_1_1320 (.ZN (n_6_1_697), .A1 (n_6_705), .A2 (n_6_1_729), .B1 (n_6_737)
    , .B2 (n_6_1_730), .C1 (n_6_2574), .C2 (n_6_1_728));
INV_X2 i_6_1_1319 (.ZN (n_6_2542), .A (n_6_1_697));
AOI222_X1 i_6_1_1318 (.ZN (n_6_1_696), .A1 (n_6_704), .A2 (n_6_1_729), .B1 (n_6_736)
    , .B2 (n_6_1_730), .C1 (n_6_2573), .C2 (n_6_1_728));
INV_X1 i_6_1_1317 (.ZN (n_6_2541), .A (n_6_1_696));
NOR2_X4 i_6_1_1316 (.ZN (sgo__n471), .A1 (n_6_1_1128), .A2 (Multiplicand[12]));
NOR2_X4 i_6_1_1315 (.ZN (sgo__n482), .A1 (Multiplicand[13]), .A2 (n_6_1_1127));
NOR2_X4 i_6_1_1314 (.ZN (n_6_1_693), .A1 (n_6_1_695), .A2 (n_6_1_694));
AND2_X1 i_6_1_1313 (.ZN (n_6_1_692), .A1 (n_6_2571), .A2 (n_6_1_693));
AOI221_X2 i_6_1_1312 (.ZN (n_6_1_691), .A (n_6_1_692), .B1 (n_6_798), .B2 (n_6_1_694)
    , .C1 (n_6_830), .C2 (n_6_1_695));
INV_X1 i_6_1_1311 (.ZN (n_6_2540), .A (n_6_1_691));
NAND2_X1 CLOCK_slo__sro_c56673 (.ZN (CLOCK_slo__sro_n51776), .A1 (slo__n28070), .A2 (n_6_1_98));
INV_X2 i_6_1_1309 (.ZN (n_6_2539), .A (n_6_1_690));
NAND2_X1 CLOCK_slo__sro_c60696 (.ZN (CLOCK_slo__sro_n55171), .A1 (n_6_2569), .A2 (n_6_1_693));
INV_X2 i_6_1_1307 (.ZN (n_6_2538), .A (CLOCK_slo__sro_n55102));
INV_X1 CLOCK_slo__sro_c61439 (.ZN (CLOCK_slo__sro_n55810), .A (n_6_2728));
INV_X2 i_6_1_1305 (.ZN (n_6_2537), .A (CLOCK_slo__sro_n55168));
NAND2_X1 slo__sro_c4826 (.ZN (slo__sro_n4618), .A1 (n_6_2085), .A2 (n_6_1_168));
INV_X2 i_6_1_1303 (.ZN (slo___n9717), .A (n_6_1_687));
INV_X2 CLOCK_slo__c69461 (.ZN (n_6_1_984), .A (CLOCK_slo__n62554));
INV_X2 i_6_1_1301 (.ZN (n_6_2535), .A (slo__sro_n8558));
AOI222_X2 i_6_1_1300 (.ZN (n_6_1_685), .A1 (n_6_824), .A2 (n_6_1_695), .B1 (n_6_792)
    , .B2 (n_6_1_694), .C1 (n_6_2566), .C2 (n_6_1_693));
INV_X2 i_6_1_1299 (.ZN (n_6_2534), .A (n_6_1_685));
NAND2_X1 slo__sro_c22563 (.ZN (slo__sro_n19570), .A1 (n_6_2320), .A2 (n_6_1_413));
INV_X2 i_6_1_1297 (.ZN (n_6_2533), .A (n_6_1_684));
NAND2_X1 slo__sro_c9322 (.ZN (slo__sro_n8685), .A1 (n_6_930), .A2 (n_6_1_625));
INV_X1 i_6_1_1295 (.ZN (n_6_2532), .A (slo__sro_n8646));
AND2_X1 slo__sro_c4419 (.ZN (slo__sro_n4245), .A1 (n_6_2724), .A2 (n_6_1_868));
INV_X1 i_6_1_1293 (.ZN (n_6_2531), .A (n_6_1_682));
NAND2_X1 CLOCK_slo__sro_c58615 (.ZN (CLOCK_slo__sro_n53420), .A1 (slo___n23359), .A2 (n_6_1244));
INV_X2 i_6_1_1291 (.ZN (n_6_2530), .A (slo__sro_n34620));
INV_X1 CLOCK_slo__c60109 (.ZN (CLOCK_slo__n54674), .A (slo__sro_n12923));
INV_X2 i_6_1_1289 (.ZN (n_6_2529), .A (CLOCK_slo__sro_n54551));
AND2_X1 CLOCK_slo__sro_c69203 (.ZN (CLOCK_slo__sro_n62332), .A1 (n_6_1401), .A2 (n_6_1_380));
INV_X1 i_6_1_1287 (.ZN (n_6_2528), .A (slo__sro_n21632));
NAND2_X1 slo__sro_c8438 (.ZN (slo__sro_n7913), .A1 (slo___n19273), .A2 (n_6_1_798));
INV_X1 i_6_1_1285 (.ZN (n_6_2527), .A (slo__sro_n7852));
NAND2_X1 slo__sro_c11066 (.ZN (slo__sro_n10273), .A1 (n_6_2645), .A2 (n_6_1_798));
INV_X1 i_6_1_1283 (.ZN (n_6_2526), .A (slo__sro_n30017));
AOI222_X2 i_6_1_1282 (.ZN (n_6_1_676), .A1 (n_6_815), .A2 (n_6_1_695), .B1 (n_6_783)
    , .B2 (n_6_1_694), .C1 (n_6_2557), .C2 (n_6_1_693));
INV_X1 i_6_1_1281 (.ZN (n_6_2525), .A (n_6_1_676));
INV_X1 CLOCK_slo__sro_c55121 (.ZN (CLOCK_slo__sro_n50403), .A (slo__sro_n35419));
INV_X1 i_6_1_1279 (.ZN (n_6_2524), .A (n_6_1_675));
NAND2_X1 slo__sro_c7881 (.ZN (slo__sro_n7408), .A1 (CLOCK_opt_ipo_n46005), .A2 (n_6_1_553));
INV_X2 i_6_1_1277 (.ZN (n_6_2523), .A (slo__sro_n7395));
INV_X2 slo__c41441 (.ZN (slo__n37528), .A (n_6_1_438));
INV_X1 i_6_1_1275 (.ZN (slo___n17357), .A (slo__sro_n7617));
AOI22_X2 slo__mro_c36955 (.ZN (slo__mro_n33300), .A1 (n_6_1948), .A2 (n_6_1_64), .B1 (n_6_2012), .B2 (n_6_1_63));
BUF_X32 drc_ipo_c29985 (.Z (drc_ipo_n26613), .A (Multiplier[18]));
NAND2_X1 CLOCK_slo__sro_c72471 (.ZN (CLOCK_slo__sro_n65089), .A1 (CLOCK_slo__sro_n65090), .A2 (CLOCK_slo__sro_n65091));
INV_X1 i_6_1_1271 (.ZN (n_6_2520), .A (slo__sro_n33788));
AOI222_X1 i_6_1_1270 (.ZN (n_6_1_670), .A1 (n_6_777), .A2 (n_6_1_694), .B1 (n_6_809)
    , .B2 (n_6_1_695), .C1 (n_6_2551), .C2 (n_6_1_693));
INV_X1 i_6_1_1269 (.ZN (n_6_2519), .A (n_6_1_670));
AOI222_X2 i_6_1_1268 (.ZN (n_6_1_669), .A1 (n_6_776), .A2 (n_6_1_694), .B1 (n_6_808)
    , .B2 (n_6_1_695), .C1 (slo___n17474), .C2 (n_6_1_693));
INV_X1 i_6_1_1267 (.ZN (n_6_2518), .A (n_6_1_669));
NAND2_X1 slo__sro_c40765 (.ZN (slo__sro_n36944), .A1 (slo__sro_n36945), .A2 (slo__sro_n36946));
INV_X1 i_6_1_1265 (.ZN (n_6_2517), .A (slo__sro_n36849));
AOI222_X2 i_6_1_1264 (.ZN (n_6_1_667), .A1 (n_6_774), .A2 (n_6_1_694), .B1 (n_6_806)
    , .B2 (n_6_1_695), .C1 (n_6_2548), .C2 (n_6_1_693));
INV_X2 i_6_1_1263 (.ZN (slo___n6972), .A (n_6_1_667));
AOI222_X2 slo__sro_c9815 (.ZN (slo__sro_n9138), .A1 (n_6_1230), .A2 (slo___n23359)
    , .B1 (n_6_1262), .B2 (slo___n23274), .C1 (n_6_2339), .C2 (n_6_1_448));
INV_X2 i_6_1_1261 (.ZN (CLOCK_slo___n52225), .A (slo__sro_n9085));
INV_X1 slo__c19332 (.ZN (slo__n17088), .A (slo__sro_n5945));
INV_X1 i_6_1_1259 (.ZN (n_6_2514), .A (slo__sro_n17074));
NAND2_X1 slo__sro_c9643 (.ZN (slo__sro_n8979), .A1 (n_6_2785), .A2 (CLOCK_sgo__n46937));
INV_X2 i_6_1_1257 (.ZN (n_6_2513), .A (slo__sro_n8916));
AOI222_X2 slo__sro_c8114 (.ZN (slo__sro_n7617), .A1 (n_6_780), .A2 (n_6_1_694), .B1 (n_6_812)
    , .B2 (n_6_1_695), .C1 (n_6_2554), .C2 (n_6_1_693));
NAND2_X1 slo__sro_c34811 (.ZN (slo__sro_n31220), .A1 (n_6_2384), .A2 (n_6_1_483));
INV_X2 i_6_1_1253 (.ZN (n_6_2511), .A (CLOCK_slo__sro_n49382));
AOI222_X1 i_6_1_1252 (.ZN (n_6_1_661), .A1 (n_6_768), .A2 (n_6_1_694), .B1 (n_6_800)
    , .B2 (n_6_1_695), .C1 (n_6_2542), .C2 (n_6_1_693));
INV_X1 i_6_1_1251 (.ZN (n_6_2510), .A (n_6_1_661));
NOR2_X4 i_6_1_1250 (.ZN (n_6_1_660), .A1 (n_6_1_1129), .A2 (Multiplicand[13]));
NOR2_X4 i_6_1_1249 (.ZN (n_6_1_659), .A1 (Multiplicand[14]), .A2 (n_6_1_1128));
NOR2_X4 i_6_1_1248 (.ZN (n_6_1_658), .A1 (slo___n23451), .A2 (slo___n23463));
AND2_X1 i_6_1_1247 (.ZN (n_6_1_657), .A1 (n_6_2540), .A2 (n_6_1_658));
AOI221_X1 i_6_1_1246 (.ZN (n_6_1_656), .A (n_6_1_657), .B1 (n_6_862), .B2 (slo___n23463)
    , .C1 (n_6_894), .C2 (slo___n23451));
INV_X1 i_6_1_1245 (.ZN (n_6_2509), .A (n_6_1_656));
AOI221_X1 i_6_1_1244 (.ZN (n_6_1_655), .A (n_6_1_657), .B1 (n_6_861), .B2 (slo___n23463)
    , .C1 (n_6_893), .C2 (slo___n23451));
INV_X1 i_6_1_1243 (.ZN (n_6_2508), .A (n_6_1_655));
CLKBUF_X1 spw__L1_c1_c76090 (.Z (n_6_2572), .A (spw__n67889));
INV_X1 i_6_1_1241 (.ZN (n_6_2507), .A (CLOCK_slo__sro_n64272));
AOI222_X2 slo__sro_c13739 (.ZN (slo__sro_n12534), .A1 (n_6_1546), .A2 (n_6_1_274)
    , .B1 (n_6_1578), .B2 (slo___n23244), .C1 (n_6_2180), .C2 (n_6_1_273));
INV_X4 i_6_1_1239 (.ZN (n_6_2506), .A (CLOCK_slo__sro_n50300));
AOI222_X2 i_6_1_1238 (.ZN (n_6_1_652), .A1 (n_6_890), .A2 (slo___n23451), .B1 (n_6_858)
    , .B2 (slo___n23463), .C1 (n_6_2537), .C2 (n_6_1_658));
INV_X2 i_6_1_1237 (.ZN (n_6_2505), .A (n_6_1_652));
AOI21_X4 slo__sro_c8218 (.ZN (slo__sro_n7705), .A (slo__mro_n33030), .B1 (n_6_750), .B2 (n_6_1_730));
INV_X1 i_6_1_1235 (.ZN (n_6_2504), .A (slo__sro_n7515));
INV_X1 slo__sro_c40637 (.ZN (slo__sro_n36837), .A (slo__sro_n17753));
INV_X2 i_6_1_1233 (.ZN (n_6_2503), .A (n_6_1_650));
AOI222_X2 i_6_1_1232 (.ZN (n_6_1_649), .A1 (n_6_887), .A2 (slo___n23451), .B1 (n_6_855)
    , .B2 (slo___n23463), .C1 (n_6_2534), .C2 (n_6_1_658));
INV_X1 i_6_1_1231 (.ZN (n_6_2502), .A (n_6_1_649));
NAND2_X1 slo__sro_c9418 (.ZN (slo__sro_n8766), .A1 (n_6_2684), .A2 (CLOCK_sgo__n46922));
INV_X2 i_6_1_1229 (.ZN (n_6_2501), .A (n_6_1_648));
INV_X2 CLOCK_slo__c71911 (.ZN (CLOCK_slo__n64621), .A (n_6_1_419));
INV_X2 i_6_1_1227 (.ZN (n_6_2500), .A (slo__sro_n32484));
NAND2_X1 slo__sro_c23579 (.ZN (slo__sro_n20509), .A1 (n_6_2127), .A2 (n_6_1_203));
INV_X1 i_6_1_1225 (.ZN (n_6_2499), .A (n_6_1_646));
INV_X1 slo__sro_c26073 (.ZN (slo__sro_n22782), .A (slo__sro_n11784));
INV_X2 i_6_1_1223 (.ZN (n_6_2498), .A (n_6_1_645));
AOI222_X2 i_6_1_1222 (.ZN (n_6_1_644), .A1 (n_6_882), .A2 (slo___n23451), .B1 (n_6_850)
    , .B2 (slo___n23463), .C1 (n_6_2529), .C2 (n_6_1_658));
INV_X2 i_6_1_1221 (.ZN (n_6_2497), .A (n_6_1_644));
NAND2_X2 slo__sro_c24582 (.ZN (slo__sro_n21438), .A1 (n_6_1433), .A2 (slo___n23229));
INV_X2 i_6_1_1219 (.ZN (n_6_2496), .A (slo__sro_n21346));
INV_X1 slo__sro_c42888 (.ZN (slo__sro_n38761), .A (slo__sro_n14590));
INV_X2 i_6_1_1217 (.ZN (n_6_2495), .A (slo__sro_n38744));
INV_X2 opt_ipo_c48207 (.ZN (opt_ipo_n43864), .A (n_0_62));
INV_X4 i_6_1_1215 (.ZN (n_6_2494), .A (slo__sro_n38758));
NAND2_X1 CLOCK_slo__sro_c69769 (.ZN (CLOCK_slo__sro_n62843), .A1 (n_6_2800), .A2 (n_6_1_973));
INV_X1 i_6_1_1213 (.ZN (n_6_2493), .A (CLOCK_slo__sro_n62783));
AOI222_X2 i_6_1_1212 (.ZN (n_6_1_639), .A1 (n_6_877), .A2 (n_6_1_660), .B1 (n_6_845)
    , .B2 (slo___n23463), .C1 (n_6_2524), .C2 (n_6_1_658));
INV_X2 i_6_1_1211 (.ZN (n_6_2492), .A (n_6_1_639));
AND2_X1 slo__sro_c36413 (.ZN (slo__sro_n32717), .A1 (n_6_2553), .A2 (n_6_1_693));
INV_X2 i_6_1_1209 (.ZN (n_6_2491), .A (slo__sro_n4338));
NOR2_X1 slo__sro_c38261 (.ZN (slo__sro_n34621), .A1 (slo__sro_n34623), .A2 (slo__sro_n34622));
INV_X1 i_6_1_1207 (.ZN (n_6_2490), .A (slo__sro_n34095));
NAND2_X1 CLOCK_slo__sro_c56071 (.ZN (CLOCK_slo__sro_n51261), .A1 (n_6_603), .A2 (n_6_1_799));
INV_X1 i_6_1_1205 (.ZN (n_6_2489), .A (slo__sro_n7557));
INV_X1 slo__sro_c41187 (.ZN (slo__sro_n37308), .A (slo__sro_n13522));
INV_X2 i_6_1_1203 (.ZN (n_6_2488), .A (n_6_1_635));
AOI222_X2 i_6_1_1202 (.ZN (n_6_1_634), .A1 (n_6_840), .A2 (slo___n23463), .B1 (n_6_872)
    , .B2 (n_6_1_660), .C1 (n_6_2519), .C2 (n_6_1_658));
INV_X2 i_6_1_1201 (.ZN (n_6_2487), .A (n_6_1_634));
INV_X1 CLOCK_sgo__sro_c51422 (.ZN (CLOCK_sgo__sro_n47200), .A (slo__sro_n7933));
INV_X2 i_6_1_1199 (.ZN (n_6_2486), .A (CLOCK_slo__sro_n59842));
INV_X1 i_6_1_1197 (.ZN (n_6_2485), .A (n_6_1_632));
NAND2_X1 slo__sro_c9795 (.ZN (slo__sro_n9124), .A1 (n_6_2278), .A2 (n_6_1_378));
INV_X2 i_6_1_1195 (.ZN (n_6_2484), .A (slo__sro_n9075));
NAND2_X1 CLOCK_slo__sro_c57659 (.ZN (CLOCK_slo__sro_n52569), .A1 (CLOCK_slo__sro_n52571), .A2 (CLOCK_slo__sro_n52570));
INV_X1 i_6_1_1193 (.ZN (n_6_2483), .A (n_6_1_630));
NAND2_X1 CLOCK_slo__sro_c54925 (.ZN (CLOCK_slo__sro_n50227), .A1 (n_6_2217), .A2 (n_6_1_308));
INV_X2 i_6_1_1191 (.ZN (n_6_2482), .A (n_6_1_629));
INV_X1 slo__sro_c24791 (.ZN (slo__sro_n21635), .A (slo__sro_n9165));
INV_X1 i_6_1_1189 (.ZN (n_6_2481), .A (slo__sro_n21560));
NAND2_X1 CLOCK_slo__sro_c69711 (.ZN (CLOCK_slo__sro_n62786), .A1 (n_6_2525), .A2 (n_6_1_658));
INV_X1 i_6_1_1187 (.ZN (n_6_2480), .A (n_6_1_627));
AOI222_X1 i_6_1_1186 (.ZN (n_6_1_626), .A1 (n_6_832), .A2 (slo___n23463), .B1 (n_6_864)
    , .B2 (n_6_1_660), .C1 (n_6_2511), .C2 (n_6_1_658));
INV_X1 i_6_1_1185 (.ZN (n_6_2479), .A (n_6_1_626));
NOR2_X1 i_6_1_1184 (.ZN (slo__n23424), .A1 (n_6_1_1130), .A2 (Multiplicand[14]));
NOR2_X4 i_6_1_1183 (.ZN (n_6_1_624), .A1 (Multiplicand[15]), .A2 (n_6_1_1129));
NOR2_X4 i_6_1_1182 (.ZN (n_6_1_623), .A1 (n_6_1_625), .A2 (slo___n23367));
AND2_X1 i_6_1_1181 (.ZN (n_6_1_622), .A1 (n_6_2509), .A2 (n_6_1_623));
AOI221_X2 i_6_1_1180 (.ZN (n_6_1_621), .A (n_6_1_622), .B1 (n_6_926), .B2 (slo___n23367)
    , .C1 (n_6_958), .C2 (n_6_1_625));
INV_X2 i_6_1_1179 (.ZN (n_6_2478), .A (n_6_1_621));
AOI221_X2 i_6_1_1178 (.ZN (n_6_1_620), .A (n_6_1_622), .B1 (n_6_925), .B2 (slo___n23367)
    , .C1 (n_6_957), .C2 (n_6_1_625));
INV_X1 i_6_1_1177 (.ZN (n_6_2477), .A (n_6_1_620));
NAND2_X1 slo__sro_c24027 (.ZN (slo__sro_n20924), .A1 (CLOCK_sgo__n46945), .A2 (opt_ipo_n24784));
INV_X2 i_6_1_1175 (.ZN (n_6_2476), .A (slo__sro_n20885));
NAND2_X2 slo__sro_c7658 (.ZN (slo__sro_n7187), .A1 (slo__sro_n7188), .A2 (slo__sro_n7189));
INV_X2 i_6_1_1173 (.ZN (n_6_2475), .A (slo__sro_n7017));
INV_X1 slo__sro_c13703 (.ZN (slo__sro_n12508), .A (n_6_2538));
INV_X2 i_6_1_1171 (.ZN (n_6_2474), .A (slo__sro_n12490));
AOI222_X2 i_6_1_1170 (.ZN (n_6_1_616), .A1 (n_6_953), .A2 (n_6_1_625), .B1 (n_6_921)
    , .B2 (slo___n23367), .C1 (n_6_2505), .C2 (n_6_1_623));
AOI222_X2 slo__sro_c6208 (.ZN (slo__sro_n5865), .A1 (n_6_1218), .A2 (slo___n23359)
    , .B1 (n_6_1250), .B2 (slo___n23274), .C1 (opt_ipo_n24251), .C2 (n_6_1_448));
INV_X1 i_6_1_1167 (.ZN (n_6_2472), .A (slo__sro_n5855));
INV_X1 CLOCK_slo__sro_c56401 (.ZN (CLOCK_slo__sro_n51544), .A (slo__sro_n36417));
INV_X2 i_6_1_1165 (.ZN (n_6_2471), .A (CLOCK_slo__sro_n51511));
AOI222_X2 i_6_1_1164 (.ZN (n_6_1_613), .A1 (n_6_950), .A2 (n_6_1_625), .B1 (n_6_918)
    , .B2 (slo___n23367), .C1 (n_6_2502), .C2 (n_6_1_623));
INV_X2 i_6_1_1163 (.ZN (n_6_2470), .A (n_6_1_613));
INV_X1 slo__sro_c32722 (.ZN (slo__sro_n29228), .A (n_6_2209));
INV_X2 i_6_1_1161 (.ZN (n_6_2469), .A (slo__sro_n19727));
AND2_X1 CLOCK_slo__sro_c55480 (.ZN (CLOCK_slo__sro_n50731), .A1 (n_6_1589), .A2 (slo___n23244));
INV_X2 i_6_1_1159 (.ZN (n_6_2468), .A (n_6_1_611));
INV_X1 CLOCK_slo__sro_c56361 (.ZN (CLOCK_slo__sro_n51512), .A (CLOCK_slo__sro_n51513));
INV_X1 i_6_1_1157 (.ZN (n_6_2467), .A (CLOCK_slo__sro_n51439));
AOI21_X1 CLOCK_slo__sro_c69752 (.ZN (CLOCK_slo__sro_n62824), .A (slo__sro_n14915)
    , .B1 (n_6_683), .B2 (n_6_1_765));
INV_X2 i_6_1_1155 (.ZN (n_6_2466), .A (CLOCK_slo__sro_n59342));
INV_X1 slo__c15705 (.ZN (slo__n14148), .A (slo__sro_n32138));
INV_X2 i_6_1_1153 (.ZN (n_6_2465), .A (slo__sro_n29443));
AND2_X1 slo__sro_c5941 (.ZN (slo__sro_n5630), .A1 (opt_ipo_n43935), .A2 (n_6_1_448));
INV_X1 i_6_1_1151 (.ZN (n_6_2464), .A (slo__sro_n20259));
AOI222_X2 slo__sro_c8183 (.ZN (n_6_1_364), .A1 (n_6_1394), .A2 (n_6_1_380), .B1 (n_6_1362)
    , .B2 (n_6_1_379), .C1 (slo__n37502), .C2 (n_6_1_378));
INV_X1 i_6_1_1149 (.ZN (n_6_2463), .A (CLOCK_slo__sro_n55687));
AND2_X1 slo__sro_c32139 (.ZN (slo__sro_n28681), .A1 (n_6_2157), .A2 (n_6_1_238));
INV_X2 i_6_1_1147 (.ZN (n_6_2462), .A (slo__sro_n28591));
AOI222_X1 i_6_1_1146 (.ZN (spw__n67656), .A1 (n_6_941), .A2 (n_6_1_625), .B1 (n_6_909)
    , .B2 (slo___n23367), .C1 (n_6_2493), .C2 (n_6_1_623));
INV_X2 i_6_1_1145 (.ZN (n_6_2461), .A (n_6_1_604));
NAND2_X1 slo__sro_c40223 (.ZN (slo__sro_n36478), .A1 (n_6_1032), .A2 (slo___n23353));
INV_X1 i_6_1_1143 (.ZN (n_6_2460), .A (CLOCK_slo__sro_n51541));
AOI222_X2 i_6_1_1142 (.ZN (n_6_1_602), .A1 (n_6_939), .A2 (n_6_1_625), .B1 (n_6_907)
    , .B2 (slo___n23367), .C1 (n_6_2491), .C2 (n_6_1_623));
INV_X2 i_6_1_1141 (.ZN (n_6_2459), .A (n_6_1_602));
INV_X8 CLOCK_slo__c53718 (.ZN (CLOCK_slo__n49141), .A (CLOCK_slo__n49140));
NAND2_X1 CLOCK_slo__sro_c54417 (.ZN (CLOCK_slo__sro_n49774), .A1 (n_6_1160), .A2 (slo___n23364));
AOI222_X2 i_6_1_1138 (.ZN (n_6_1_600), .A1 (n_6_937), .A2 (n_6_1_625), .B1 (n_6_905)
    , .B2 (slo___n23367), .C1 (n_6_2489), .C2 (n_6_1_623));
INV_X2 i_6_1_1137 (.ZN (n_6_2457), .A (n_6_1_600));
NAND2_X1 CLOCK_slo__sro_c55401 (.ZN (CLOCK_slo__sro_n50659), .A1 (n_6_1070), .A2 (slo___n23457));
INV_X2 i_6_1_1135 (.ZN (n_6_2456), .A (CLOCK_slo__sro_n50608));
AND2_X1 slo__sro_c6377 (.ZN (slo__sro_n6021), .A1 (n_6_2317), .A2 (n_6_1_413));
INV_X2 i_6_1_1133 (.ZN (n_6_2455), .A (slo__sro_n31559));
INV_X1 slo__sro_c23687 (.ZN (slo__sro_n20614), .A (CLOCK_sgo__n46950));
INV_X2 i_6_1_1131 (.ZN (slo___n17886), .A (slo__sro_n42341));
NAND2_X1 slo__sro_c24841 (.ZN (slo__sro_n21678), .A1 (n_6_1_734), .A2 (n_6_1_728));
INV_X1 i_6_1_1129 (.ZN (n_6_2453), .A (slo__sro_n21662));
AOI222_X2 slo__sro_c41045 (.ZN (slo__sro_n37192), .A1 (n_6_680), .A2 (n_6_1_765), .B1 (n_6_648)
    , .B2 (n_6_1_764), .C1 (n_6_2612), .C2 (n_6_1_763));
INV_X2 i_6_1_1127 (.ZN (n_6_2452), .A (n_6_1_595));
NAND2_X1 slo__sro_c7946 (.ZN (slo__sro_n7465), .A1 (slo__sro_n7466), .A2 (slo__sro_n7467));
INV_X1 i_6_1_1125 (.ZN (n_6_2451), .A (slo__sro_n32044));
AND2_X1 slo__sro_c9389 (.ZN (slo__sro_n8742), .A1 (n_6_2721), .A2 (n_6_1_868));
INV_X2 i_6_1_1123 (.ZN (n_6_2450), .A (n_6_1_593));
AOI222_X2 i_6_1_1122 (.ZN (n_6_1_592), .A1 (n_6_897), .A2 (slo___n23367), .B1 (n_6_929)
    , .B2 (n_6_1_625), .C1 (n_6_2481), .C2 (n_6_1_623));
INV_X2 i_6_1_1121 (.ZN (slo__n31336), .A (n_6_1_592));
AOI222_X2 i_6_1_1120 (.ZN (n_6_1_591), .A1 (n_6_896), .A2 (slo___n23367), .B1 (n_6_928)
    , .B2 (n_6_1_625), .C1 (n_6_2480), .C2 (n_6_1_623));
INV_X2 i_6_1_1119 (.ZN (n_6_2448), .A (n_6_1_591));
NOR2_X4 i_6_1_1118 (.ZN (n_6_1_590), .A1 (n_6_1_1131), .A2 (Multiplicand[15]));
NOR2_X4 i_6_1_1117 (.ZN (n_6_1_589), .A1 (Multiplicand[16]), .A2 (n_6_1_1130));
NOR2_X4 i_6_1_1116 (.ZN (n_6_1_588), .A1 (slo___n23218), .A2 (slo___n23232));
AND2_X1 i_6_1_1115 (.ZN (n_6_1_587), .A1 (n_6_2478), .A2 (n_6_1_588));
AOI221_X2 i_6_1_1114 (.ZN (n_6_1_586), .A (n_6_1_587), .B1 (n_6_990), .B2 (slo___n23232)
    , .C1 (n_6_1022), .C2 (slo___n23218));
INV_X2 i_6_1_1113 (.ZN (n_6_2447), .A (n_6_1_586));
AOI21_X1 CLOCK_slo__sro_c56906 (.ZN (CLOCK_slo__sro_n51958), .A (slo__sro_n12328)
    , .B1 (n_6_364), .B2 (n_6_1_940));
INV_X4 i_6_1_1111 (.ZN (n_6_2446), .A (n_6_1_585));
AND2_X1 slo__sro_c25707 (.ZN (slo__sro_n22458), .A1 (n_6_2236), .A2 (n_6_1_343));
CLKBUF_X1 CLOCK_slo___L1_c1_c57283 (.Z (slo___n16283), .A (CLOCK_slo___n52225));
NAND2_X1 slo__sro_c37467 (.ZN (slo__sro_n33790), .A1 (n_6_2552), .A2 (n_6_1_693));
INV_X2 i_6_1_1107 (.ZN (n_6_2444), .A (slo__sro_n33776));
NAND2_X1 slo__sro_c8813 (.ZN (slo__sro_n8245), .A1 (n_6_2766), .A2 (CLOCK_sgo__n46937));
AND2_X1 slo__sro_c32943 (.ZN (slo__sro_n29444), .A1 (n_6_945), .A2 (n_6_1_625));
AOI222_X2 i_6_1_1104 (.ZN (n_6_1_581), .A1 (n_6_1017), .A2 (slo___n23218), .B1 (n_6_985)
    , .B2 (slo___n23232), .C1 (n_6_2474), .C2 (n_6_1_588));
INV_X2 i_6_1_1103 (.ZN (n_6_2442), .A (n_6_1_581));
NAND2_X1 slo__sro_c42474 (.ZN (slo__sro_n38411), .A1 (n_6_2234), .A2 (n_6_1_343));
INV_X2 slo__c42215 (.ZN (slo__n38193), .A (slo__sro_n20680));
AOI221_X2 slo__sro_c37457 (.ZN (slo__sro_n33776), .A (slo__sro_n33777), .B1 (n_6_987)
    , .B2 (slo___n23232), .C1 (n_6_1019), .C2 (slo___n23218));
INV_X1 i_6_1_1099 (.ZN (n_6_2440), .A (slo__sro_n33466));
AOI222_X2 slo__sro_c37135 (.ZN (slo__sro_n33466), .A1 (n_6_1015), .A2 (slo___n23218)
    , .B1 (n_6_983), .B2 (slo___n23232), .C1 (n_6_2472), .C2 (n_6_1_588));
INV_X2 i_6_1_1097 (.ZN (n_6_2439), .A (slo__sro_n33384));
INV_X1 CLOCK_opt_ipo_c50073 (.ZN (CLOCK_opt_ipo_n45730), .A (n_6_1_58));
INV_X1 i_6_1_1095 (.ZN (n_6_2438), .A (n_6_1_577));
NAND2_X1 CLOCK_slo__sro_c66052 (.ZN (CLOCK_slo__sro_n59535), .A1 (n_6_2094), .A2 (n_6_1_168));
INV_X2 i_6_1_1093 (.ZN (n_6_2437), .A (slo__sro_n6088));
AOI222_X2 i_6_1_1092 (.ZN (n_6_1_575), .A1 (n_6_1011), .A2 (slo___n23218), .B1 (n_6_979)
    , .B2 (slo___n23232), .C1 (n_6_2468), .C2 (n_6_1_588));
INV_X1 i_6_1_1091 (.ZN (n_6_2436), .A (n_6_1_575));
AOI21_X4 slo__sro_c10487 (.ZN (slo__sro_n9753), .A (slo__sro_n9754), .B1 (n_6_1463), .B2 (n_6_1_345));
INV_X1 i_6_1_1089 (.ZN (n_6_2435), .A (n_6_1_574));
NAND2_X1 slo__sro_c33834 (.ZN (slo__sro_n30285), .A1 (slo__sro_n30286), .A2 (slo__sro_n30287));
NAND2_X1 slo__sro_c44140 (.ZN (Product[60]), .A1 (slo__sro_n39768), .A2 (slo__sro_n39769));
INV_X2 i_6_1_1085 (.ZN (n_6_2433), .A (n_6_1_572));
AOI222_X2 i_6_1_1084 (.ZN (n_6_1_571), .A1 (n_6_1007), .A2 (slo___n23218), .B1 (n_6_975)
    , .B2 (slo___n23232), .C1 (n_6_2464), .C2 (n_6_1_588));
INV_X2 i_6_1_1083 (.ZN (n_6_2432), .A (n_6_1_571));
INV_X1 slo__mro_c36717 (.ZN (slo__mro_n33047), .A (n_6_1_834));
INV_X2 i_6_1_1081 (.ZN (n_6_2431), .A (slo__sro_n7689));
INV_X1 slo__sro_c23024 (.ZN (slo__sro_n19999), .A (n_6_1_448));
INV_X2 i_6_1_1079 (.ZN (n_6_2430), .A (slo__sro_n19958));
INV_X1 slo__sro_c23023 (.ZN (slo__sro_n20000), .A (n_6_2335));
INV_X1 i_6_1_1077 (.ZN (n_6_2429), .A (slo__sro_n19970));
NAND2_X1 CLOCK_slo__sro_c54832 (.ZN (CLOCK_slo__sro_n50141), .A1 (n_6_2284), .A2 (n_6_1_378));
INV_X4 CLOCK_slo__c53453 (.ZN (n_6_1_150), .A (CLOCK_slo__n48906));
NAND2_X1 slo__sro_c42376 (.ZN (slo__sro_n38324), .A1 (n_6_1_273), .A2 (n_6_2182));
INV_X1 slo__sro_c40160 (.ZN (slo__sro_n36418), .A (n_6_1_623));
NAND2_X1 slo__sro_c31434 (.ZN (slo__sro_n28008), .A1 (n_6_2559), .A2 (n_6_1_693));
INV_X1 i_6_1_1071 (.ZN (n_6_2426), .A (CLOCK_slo__sro_n52136));
INV_X1 i_6_1_1069 (.ZN (n_6_2425), .A (slo__sro_n28419));
AOI221_X2 slo__sro_c45412 (.ZN (slo__sro_n40936), .A (slo__sro_n40937), .B1 (n_6_1227)
    , .B2 (slo___n23359), .C1 (n_6_1259), .C2 (slo___n23274));
INV_X1 i_6_1_1067 (.ZN (n_6_2424), .A (n_6_1_563));
CLKBUF_X1 slo___L1_c1_c20702 (.Z (n_6_2099), .A (CLOCK_slo__n56418));
INV_X4 i_6_1_1065 (.ZN (n_6_2423), .A (n_6_1_562));
BUF_X1 spc__L1_c74527 (.Z (spc__n66318), .A (n_6_1_134));
INV_X1 i_6_1_1063 (.ZN (n_6_2422), .A (CLOCK_slo__sro_n51132));
AND2_X1 slo__sro_c7911 (.ZN (slo__sro_n7436), .A1 (n_6_2394), .A2 (n_6_1_518));
INV_X2 i_6_1_1061 (.ZN (n_6_2421), .A (slo__sro_n41029));
AOI222_X2 slo__sro_c7740 (.ZN (slo__sro_n7270), .A1 (n_6_994), .A2 (slo___n23218)
    , .B1 (n_6_962), .B2 (slo___n23232), .C1 (n_6_2451), .C2 (n_6_1_588));
INV_X2 i_6_1_1059 (.ZN (n_6_2420), .A (slo__sro_n7186));
NAND2_X1 slo__sro_c7776 (.ZN (slo__sro_n7309), .A1 (n_6_2280), .A2 (n_6_1_378));
INV_X2 i_6_1_1057 (.ZN (n_6_2419), .A (slo__sro_n7270));
INV_X1 CLOCK_slo__sro_c60518 (.ZN (CLOCK_slo__sro_n55021), .A (slo___n23359));
INV_X2 i_6_1_1055 (.ZN (n_6_2418), .A (n_6_1_557));
AOI222_X1 i_6_1_1054 (.ZN (n_6_1_556), .A1 (n_6_960), .A2 (slo___n23232), .B1 (n_6_992)
    , .B2 (slo___n23218), .C1 (slo__n31336), .C2 (n_6_1_588));
INV_X1 i_6_1_1053 (.ZN (n_6_2417), .A (n_6_1_556));
NOR2_X4 i_6_1_1052 (.ZN (n_6_1_555), .A1 (n_6_1_1132), .A2 (Multiplicand[16]));
NOR2_X1 i_6_1_1051 (.ZN (slo__n41748), .A1 (Multiplicand[17]), .A2 (n_6_1_1131));
NOR2_X4 i_6_1_1050 (.ZN (n_6_1_553), .A1 (slo___n23457), .A2 (n_6_1_554));
AND2_X1 i_6_1_1049 (.ZN (n_6_1_552), .A1 (n_6_2447), .A2 (n_6_1_553));
AOI21_X2 slo__sro_c40766 (.ZN (n_6_1_595), .A (slo__sro_n36944), .B1 (n_6_900), .B2 (slo___n23367));
INV_X1 i_6_1_1047 (.ZN (n_6_2416), .A (slo__sro_n36810));
AOI221_X1 i_6_1_1046 (.ZN (n_6_1_550), .A (n_6_1_552), .B1 (n_6_1053), .B2 (n_6_1_554)
    , .C1 (n_6_1085), .C2 (slo___n23457));
INV_X1 i_6_1_1045 (.ZN (n_6_2415), .A (n_6_1_550));
NAND2_X1 CLOCK_slo__sro_c65773 (.ZN (CLOCK_slo__sro_n59283), .A1 (n_6_2835), .A2 (CLOCK_sgo__n46950));
INV_X1 i_6_1_1043 (.ZN (n_6_2414), .A (n_6_1_549));
BUF_X8 drc_ipo_c29977 (.Z (drc_ipo_n26600), .A (slo__n4958));
INV_X2 i_6_1_1041 (.ZN (n_6_2413), .A (n_6_1_548));
AOI21_X1 slo__sro_c12767 (.ZN (slo__sro_n11706), .A (slo__sro_n11707), .B1 (n_6_139), .B2 (n_6_1_1044));
INV_X2 i_6_1_1039 (.ZN (n_6_2412), .A (n_6_1_547));
NAND2_X1 slo__sro_c22813 (.ZN (slo__sro_n19807), .A1 (n_6_1_835), .A2 (n_6_561));
INV_X4 i_6_1_1037 (.ZN (n_6_2411), .A (slo__sro_n30995));
NAND2_X1 CLOCK_sgo__sro_c51748 (.ZN (CLOCK_sgo__sro_n47470), .A1 (slo__n33292), .A2 (n_6_1_168));
INV_X2 i_6_1_1035 (.ZN (n_6_2410), .A (n_6_1_545));
NAND2_X1 slo__sro_c5046 (.ZN (slo__sro_n4816), .A1 (n_6_2909), .A2 (slo__n13799));
INV_X1 i_6_1_1033 (.ZN (n_6_2409), .A (slo__sro_n4784));
AND2_X1 slo__sro_c8727 (.ZN (slo__sro_n8171), .A1 (n_6_2762), .A2 (CLOCK_sgo__n46937));
INV_X2 i_6_1_1031 (.ZN (n_6_2408), .A (slo__sro_n8092));
AOI222_X2 i_6_1_1030 (.ZN (slo__n41747), .A1 (n_6_1077), .A2 (slo___n23457), .B1 (n_6_1045)
    , .B2 (n_6_1_554), .C1 (n_6_2439), .C2 (n_6_1_553));
NAND2_X1 slo__sro_c46337 (.ZN (slo__sro_n41833), .A1 (n_6_2848), .A2 (CLOCK_sgo__n46950));
NAND2_X2 slo__sro_c35456 (.ZN (slo__sro_n31818), .A1 (n_6_389), .A2 (n_6_1_904));
INV_X2 i_6_1_1027 (.ZN (n_6_2406), .A (slo__sro_n31798));
AOI222_X2 i_6_1_1026 (.ZN (n_6_1_540), .A1 (n_6_1075), .A2 (slo___n23457), .B1 (n_6_1043)
    , .B2 (n_6_1_554), .C1 (n_6_2437), .C2 (n_6_1_553));
INV_X1 i_6_1_1025 (.ZN (n_6_2405), .A (n_6_1_540));
AOI222_X1 i_6_1_1024 (.ZN (n_6_1_539), .A1 (n_6_1074), .A2 (slo___n23457), .B1 (n_6_1042)
    , .B2 (n_6_1_554), .C1 (n_6_2436), .C2 (n_6_1_553));
INV_X1 i_6_1_1023 (.ZN (n_6_2404), .A (n_6_1_539));
NOR2_X1 CLOCK_slo__sro_c70043 (.ZN (n_6_1_849), .A1 (CLOCK_slo__sro_n51619), .A2 (CLOCK_slo__sro_n63090));
INV_X2 i_6_1_1021 (.ZN (n_6_2403), .A (CLOCK_slo__sro_n63004));
AND2_X1 CLOCK_slo__sro_c56967 (.ZN (CLOCK_slo__sro_n52005), .A1 (n_6_508), .A2 (n_6_1_870));
INV_X1 i_6_1_1019 (.ZN (n_6_2402), .A (CLOCK_slo__sro_n54053));
NAND2_X1 CLOCK_slo__sro_c55400 (.ZN (CLOCK_slo__sro_n50660), .A1 (n_6_2432), .A2 (n_6_1_553));
INV_X2 i_6_1_1017 (.ZN (n_6_2401), .A (CLOCK_slo__n65456));
AND2_X1 CLOCK_slo__sro_c53654 (.ZN (CLOCK_slo__sro_n49084), .A1 (slo___n17155), .A2 (n_6_1_448));
INV_X1 i_6_1_1015 (.ZN (slo___n15030), .A (CLOCK_slo__sro_n50657));
AOI222_X2 i_6_1_1014 (.ZN (slo__n35115), .A1 (n_6_1069), .A2 (slo___n23457), .B1 (n_6_1037)
    , .B2 (n_6_1_554), .C1 (n_6_2431), .C2 (n_6_1_553));
NAND2_X1 slo__sro_c38840 (.ZN (slo__sro_n35185), .A1 (n_6_661), .A2 (n_6_1_764));
NAND2_X1 slo__sro_c8352 (.ZN (slo__sro_n7834), .A1 (n_6_123), .A2 (n_6_1_1080));
INV_X2 i_6_1_1011 (.ZN (n_6_2398), .A (CLOCK_slo__sro_n55059));
AOI221_X2 slo__sro_c7213 (.ZN (slo__sro_n6790), .A (slo__sro_n6791), .B1 (n_6_1326)
    , .B2 (slo___n43257), .C1 (n_6_1294), .C2 (n_6_1_414));
INV_X2 i_6_1_1009 (.ZN (n_6_2397), .A (n_6_1_532));
NAND2_X1 slo__sro_c7897 (.ZN (slo__sro_n7423), .A1 (n_6_2453), .A2 (n_6_1_588));
AND2_X1 CLOCK_slo__sro_c60559 (.ZN (CLOCK_slo__sro_n55060), .A1 (n_6_1036), .A2 (slo___n23353));
INV_X1 slo__sro_c35773 (.ZN (slo__sro_n32120), .A (n_6_2392));
INV_X4 i_6_1_1005 (.ZN (n_6_2395), .A (slo__sro_n7331));
NAND2_X1 slo__sro_c40639 (.ZN (slo__sro_n36835), .A1 (slo__sro_n36836), .A2 (slo__sro_n36837));
INV_X1 i_6_1_1003 (.ZN (n_6_2394), .A (slo__sro_n36476));
AOI222_X2 i_6_1_1002 (.ZN (n_6_1_528), .A1 (n_6_1063), .A2 (slo___n23457), .B1 (n_6_1031)
    , .B2 (slo___n23353), .C1 (n_6_2425), .C2 (n_6_1_553));
INV_X2 i_6_1_1001 (.ZN (n_6_2393), .A (n_6_1_528));
NAND2_X1 slo__sro_c8201 (.ZN (slo__sro_n7690), .A1 (slo__sro_n7691), .A2 (slo__sro_n7692));
INV_X2 i_6_1_999 (.ZN (n_6_2392), .A (slo__sro_n7633));
AOI222_X2 i_6_1_998 (.ZN (n_6_1_526), .A1 (n_6_1029), .A2 (slo___n23353), .B1 (n_6_1061)
    , .B2 (slo___n23457), .C1 (n_6_2423), .C2 (n_6_1_553));
INV_X2 i_6_1_997 (.ZN (n_6_2391), .A (n_6_1_526));
NAND2_X1 slo__sro_c7292 (.ZN (slo__sro_n6871), .A1 (n_6_1172), .A2 (slo___n23364));
INV_X2 i_6_1_995 (.ZN (n_6_2390), .A (slo__sro_n6852));
AOI222_X2 i_6_1_994 (.ZN (n_6_1_524), .A1 (n_6_1027), .A2 (slo___n23353), .B1 (n_6_1059)
    , .B2 (slo___n23457), .C1 (n_6_2421), .C2 (n_6_1_553));
INV_X2 i_6_1_993 (.ZN (slo___n6965), .A (n_6_1_524));
AOI222_X1 i_6_1_992 (.ZN (n_6_1_523), .A1 (n_6_1026), .A2 (slo___n23353), .B1 (n_6_1058)
    , .B2 (slo___n23457), .C1 (n_6_2420), .C2 (n_6_1_553));
INV_X1 CLOCK_sgo__sro_c51591 (.ZN (CLOCK_sgo__sro_n47339), .A (slo__sro_n5417));
AOI21_X2 slo__sro_c7779 (.ZN (slo__sro_n7306), .A (slo__sro_n7307), .B1 (n_6_1393), .B2 (n_6_1_380));
INV_X2 i_6_1_989 (.ZN (slo___n7115), .A (n_6_1_522));
AOI222_X1 i_6_1_988 (.ZN (n_6_1_521), .A1 (n_6_1024), .A2 (slo___n23353), .B1 (n_6_1056)
    , .B2 (slo___n23457), .C1 (n_6_2418), .C2 (n_6_1_553));
INV_X1 i_6_1_987 (.ZN (n_6_2386), .A (n_6_1_521));
NOR2_X1 i_6_1_986 (.ZN (n_6_1_520), .A1 (n_6_1_1133), .A2 (Multiplicand[17]));
NOR2_X4 i_6_1_985 (.ZN (n_6_1_519), .A1 (Multiplicand[18]), .A2 (n_6_1_1132));
NOR2_X4 i_6_1_984 (.ZN (n_6_1_518), .A1 (slo___n23268), .A2 (slo___n23277));
AND2_X1 i_6_1_983 (.ZN (n_6_1_517), .A1 (n_6_2416), .A2 (n_6_1_518));
AOI221_X1 i_6_1_982 (.ZN (n_6_1_516), .A (n_6_1_517), .B1 (n_6_1118), .B2 (slo___n23277)
    , .C1 (n_6_1150), .C2 (slo___n23268));
NAND2_X1 CLOCK_sgo__sro_c51423 (.ZN (CLOCK_sgo__sro_n47199), .A1 (n_6_356), .A2 (n_6_1_940));
AOI221_X2 i_6_1_980 (.ZN (n_6_1_515), .A (n_6_1_517), .B1 (n_6_1117), .B2 (slo___n23277)
    , .C1 (n_6_1149), .C2 (slo___n23268));
INV_X2 i_6_1_979 (.ZN (n_6_2384), .A (n_6_1_515));
AND2_X1 slo__sro_c20202 (.ZN (slo__sro_n17761), .A1 (opt_ipo_n24966), .A2 (n_6_1_553));
INV_X1 i_6_1_977 (.ZN (n_6_2383), .A (n_6_1_514));
NAND2_X1 slo__sro_c12765 (.ZN (slo__sro_n11708), .A1 (n_6_1_1045), .A2 (n_6_171));
INV_X2 i_6_1_975 (.ZN (n_6_2382), .A (n_6_1_513));
INV_X1 slo__c20144 (.ZN (slo__n17713), .A (n_6_1_124));
INV_X2 i_6_1_973 (.ZN (n_6_2381), .A (CLOCK_slo__sro_n58904));
NAND2_X1 CLOCK_slo__sro_c53955 (.ZN (CLOCK_slo__sro_n49350), .A1 (opt_ipo_n24431), .A2 (n_6_1_343));
INV_X1 i_6_1_971 (.ZN (n_6_2380), .A (n_6_1_511));
NAND2_X1 slo__sro_c31251 (.ZN (slo__sro_n27838), .A1 (n_6_2793), .A2 (n_6_1_973));
INV_X2 i_6_1_969 (.ZN (n_6_2379), .A (slo__sro_n27822));
AOI222_X2 i_6_1_968 (.ZN (n_6_1_509), .A1 (n_6_1143), .A2 (n_6_1_520), .B1 (n_6_1111)
    , .B2 (slo___n23277), .C1 (n_6_2410), .C2 (n_6_1_518));
INV_X2 i_6_1_967 (.ZN (n_6_2378), .A (n_6_1_509));
INV_X1 slo__sro_c5016 (.ZN (slo__sro_n4787), .A (opt_ipo_n24743));
INV_X1 i_6_1_965 (.ZN (n_6_2377), .A (slo__sro_n4774));
AOI222_X2 i_6_1_964 (.ZN (n_6_1_507), .A1 (n_6_1141), .A2 (slo___n23268), .B1 (n_6_1109)
    , .B2 (slo___n23277), .C1 (n_6_2408), .C2 (n_6_1_518));
INV_X1 i_6_1_963 (.ZN (n_6_2376), .A (n_6_1_507));
NAND2_X1 slo__sro_c37893 (.ZN (slo__sro_n34279), .A1 (n_6_2287), .A2 (n_6_1_378));
INV_X2 i_6_1_961 (.ZN (n_6_2375), .A (slo__sro_n34087));
NAND2_X1 slo__sro_c32860 (.ZN (slo__sro_n29365), .A1 (n_6_1_588), .A2 (n_6_2466));
INV_X1 i_6_1_959 (.ZN (n_6_2374), .A (n_6_1_505));
AOI222_X2 i_6_1_958 (.ZN (n_6_1_504), .A1 (n_6_1138), .A2 (slo___n23268), .B1 (n_6_1106)
    , .B2 (slo___n23277), .C1 (n_6_2405), .C2 (n_6_1_518));
INV_X1 i_6_1_957 (.ZN (n_6_2373), .A (n_6_1_504));
AND2_X1 slo__sro_c5166 (.ZN (slo__sro_n4923), .A1 (n_6_2252), .A2 (n_6_1_343));
INV_X1 i_6_1_955 (.ZN (n_6_2372), .A (slo__sro_n4880));
AOI222_X2 slo__sro_c6198 (.ZN (slo__sro_n5855), .A1 (n_6_952), .A2 (n_6_1_625), .B1 (n_6_920)
    , .B2 (slo___n23367), .C1 (n_6_2504), .C2 (n_6_1_623));
INV_X2 i_6_1_953 (.ZN (n_6_2371), .A (CLOCK_slo__sro_n51979));
AOI222_X2 i_6_1_952 (.ZN (n_6_1_501), .A1 (n_6_1135), .A2 (slo___n23268), .B1 (n_6_1103)
    , .B2 (slo___n23277), .C1 (n_6_2402), .C2 (n_6_1_518));
INV_X2 i_6_1_951 (.ZN (n_6_2370), .A (n_6_1_501));
NAND2_X1 slo__sro_c37895 (.ZN (slo__sro_n34277), .A1 (CLOCK_slo__mro_n63339), .A2 (slo__sro_n34279));
INV_X2 i_6_1_949 (.ZN (slo___n19058), .A (slo__sro_n33814));
AOI21_X2 slo__sro_c6221 (.ZN (slo__sro_n5875), .A (slo__sro_n5876), .B1 (n_6_1641), .B2 (drc_ipo_n26601));
INV_X2 i_6_1_947 (.ZN (n_6_2368), .A (slo__sro_n5794));
INV_X1 slo__sro_c23456 (.ZN (slo__sro_n20396), .A (n_6_2277));
INV_X1 i_6_1_945 (.ZN (n_6_2367), .A (slo__sro_n20321));
INV_X1 slo__L1_c2_c34250 (.ZN (slo__n30671), .A (slo__sro_n36913));
INV_X2 i_6_1_943 (.ZN (n_6_2366), .A (slo__sro_n30284));
AOI222_X2 i_6_1_942 (.ZN (n_6_1_496), .A1 (n_6_1130), .A2 (slo___n23268), .B1 (n_6_1098)
    , .B2 (slo___n23277), .C1 (n_6_2397), .C2 (n_6_1_518));
INV_X1 i_6_1_941 (.ZN (n_6_2365), .A (n_6_1_496));
AND2_X1 slo__sro_c10663 (.ZN (slo__sro_n9916), .A1 (n_6_2291), .A2 (n_6_1_378));
INV_X2 i_6_1_939 (.ZN (n_6_2364), .A (slo__sro_n9845));
NAND2_X1 slo__sro_c41086 (.ZN (slo__sro_n37222), .A1 (slo__sro_n37223), .A2 (slo__sro_n37224));
BUF_X32 drc_ipo_c29978 (.Z (drc_ipo_n26601), .A (n_6_1_240));
AND2_X1 slo__sro_c7923 (.ZN (slo__sro_n7448), .A1 (n_6_2717), .A2 (n_6_1_868));
INV_X1 i_6_1_935 (.ZN (n_6_2362), .A (slo__sro_n7435));
AND2_X1 slo__sro_c12503 (.ZN (slo__sro_n11483), .A1 (n_6_2748), .A2 (CLOCK_sgo__n46934));
INV_X2 i_6_1_933 (.ZN (n_6_2361), .A (n_6_1_492));
NAND2_X1 slo__sro_c34286 (.ZN (slo__sro_n30706), .A1 (n_6_1_904), .A2 (n_6_412));
INV_X2 i_6_1_931 (.ZN (n_6_2360), .A (slo__sro_n32117));
INV_X1 slo__c19655 (.ZN (slo__n17338), .A (slo__sro_n11383));
INV_X2 i_6_1_929 (.ZN (n_6_2359), .A (slo__sro_n31087));
AOI222_X2 i_6_1_928 (.ZN (n_6_1_489), .A1 (n_6_1091), .A2 (slo___n23277), .B1 (n_6_1123)
    , .B2 (slo___n23268), .C1 (n_6_2390), .C2 (n_6_1_518));
INV_X2 i_6_1_927 (.ZN (slo___n17582), .A (n_6_1_489));
INV_X1 i_6_1_925 (.ZN (n_6_2357), .A (n_6_1_488));
AOI222_X2 i_6_1_924 (.ZN (n_6_1_487), .A1 (n_6_1089), .A2 (slo___n23277), .B1 (n_6_1121)
    , .B2 (slo___n23268), .C1 (n_6_2388), .C2 (n_6_1_518));
INV_X2 i_6_1_923 (.ZN (n_6_2356), .A (n_6_1_487));
AOI222_X1 i_6_1_922 (.ZN (n_6_1_486), .A1 (n_6_1088), .A2 (slo___n23277), .B1 (n_6_1120)
    , .B2 (slo___n23268), .C1 (slo___n7115), .C2 (n_6_1_518));
INV_X1 i_6_1_921 (.ZN (n_6_2355), .A (n_6_1_486));
NOR2_X4 i_6_1_920 (.ZN (n_6_1_485), .A1 (n_6_1_1134), .A2 (Multiplicand[18]));
NOR2_X4 i_6_1_919 (.ZN (n_6_1_484), .A1 (Multiplicand[19]), .A2 (n_6_1_1133));
NOR2_X4 i_6_1_918 (.ZN (n_6_1_483), .A1 (slo___n23466), .A2 (slo___n23364));
AND2_X1 i_6_1_917 (.ZN (n_6_1_482), .A1 (opt_ipo_n45144), .A2 (n_6_1_483));
AOI221_X2 i_6_1_916 (.ZN (n_6_1_481), .A (n_6_1_482), .B1 (n_6_1182), .B2 (slo___n23364)
    , .C1 (n_6_1214), .C2 (slo___n23466));
INV_X2 i_6_1_915 (.ZN (n_6_2354), .A (n_6_1_481));
NAND2_X1 CLOCK_slo__sro_c57141 (.ZN (CLOCK_slo__sro_n52138), .A1 (n_6_1001), .A2 (slo___n23218));
NAND2_X1 CLOCK_slo__sro_c68064 (.ZN (CLOCK_slo__sro_n61297), .A1 (n_6_2883), .A2 (slo__n13799));
NAND2_X1 slo__sro_c34831 (.ZN (slo__sro_n31237), .A1 (n_6_2303), .A2 (n_6_1_413));
INV_X4 i_6_1_911 (.ZN (n_6_2352), .A (n_6_1_479));
INV_X1 slo__sro_c45410 (.ZN (slo__sro_n40938), .A (n_6_1_448));
INV_X1 i_6_1_909 (.ZN (n_6_2351), .A (CLOCK_slo__sro_n49022));
NAND2_X1 slo__sro_c42874 (.ZN (slo__sro_n38747), .A1 (n_6_2527), .A2 (n_6_1_658));
INV_X2 i_6_1_907 (.ZN (n_6_2350), .A (slo__sro_n38698));
AOI21_X2 slo__c20171 (.ZN (slo__n17737), .A (slo__sro_n7465), .B1 (n_6_1187), .B2 (slo___n23466));
INV_X1 i_6_1_905 (.ZN (n_6_2349), .A (slo__sro_n17646));
AOI222_X2 i_6_1_904 (.ZN (n_6_1_475), .A1 (n_6_1208), .A2 (slo___n23466), .B1 (n_6_1176)
    , .B2 (slo___n23364), .C1 (n_6_2380), .C2 (n_6_1_483));
INV_X2 i_6_1_903 (.ZN (n_6_2348), .A (n_6_1_475));
NAND2_X1 slo__sro_c31868 (.ZN (slo__sro_n28422), .A1 (n_6_2457), .A2 (n_6_1_588));
INV_X1 CLOCK_slo__sro_c55631 (.ZN (CLOCK_slo__sro_n50864), .A (slo__sro_n10839));
NAND2_X1 slo__sro_c22812 (.ZN (slo__sro_n19808), .A1 (n_6_2683), .A2 (CLOCK_sgo__n46922));
INV_X2 i_6_1_899 (.ZN (n_6_2346), .A (slo__sro_n19695));
NAND2_X1 slo__sro_c19676 (.ZN (slo__sro_n17353), .A1 (n_6_913), .A2 (slo___n23367));
INV_X2 i_6_1_897 (.ZN (n_6_2345), .A (slo__sro_n17330));
AOI222_X2 slo__sro_c7313 (.ZN (n_6_1_488), .A1 (n_6_1122), .A2 (slo___n23268), .B1 (n_6_1090)
    , .B2 (slo___n23277), .C1 (slo___n6965), .C2 (n_6_1_518));
INV_X2 i_6_1_895 (.ZN (n_6_2344), .A (slo__sro_n6869));
AOI222_X2 CLOCK_slo__sro_c72402 (.ZN (CLOCK_slo__sro_n65030), .A1 (n_6_193), .A2 (n_6_1_1009)
    , .B1 (n_6_225), .B2 (n_6_1_1010), .C1 (slo___n5717), .C2 (CLOCK_sgo__n46950));
INV_X1 i_6_1_893 (.ZN (n_6_2343), .A (n_6_1_470));
AOI222_X1 i_6_1_892 (.ZN (n_6_1_469), .A1 (n_6_1202), .A2 (slo___n23466), .B1 (n_6_1170)
    , .B2 (slo___n23364), .C1 (n_6_2374), .C2 (n_6_1_483));
INV_X2 i_6_1_891 (.ZN (n_6_2342), .A (n_6_1_469));
AOI222_X2 slo__sro_c37700 (.ZN (slo__sro_n34087), .A1 (n_6_1108), .A2 (slo___n23277)
    , .B1 (n_6_1140), .B2 (n_6_1_520), .C1 (n_6_1_542), .C2 (n_6_1_518));
INV_X2 i_6_1_889 (.ZN (n_6_2341), .A (slo__sro_n9805));
NAND2_X1 CLOCK_slo__sro_c57759 (.ZN (CLOCK_slo__sro_n52670), .A1 (slo___n23232), .A2 (n_6_982));
INV_X2 i_6_1_887 (.ZN (n_6_2340), .A (slo__sro_n9268));
NAND2_X1 slo__sro_c9584 (.ZN (slo__sro_n8917), .A1 (slo__sro_n8918), .A2 (slo__sro_n8919));
INV_X1 i_6_1_885 (.ZN (n_6_2339), .A (slo__sro_n8900));
INV_X1 slo__sro_c6032 (.ZN (slo__sro_n5713), .A (opt_ipo_n24861));
INV_X1 i_6_1_883 (.ZN (n_6_2338), .A (slo__sro_n5678));
AOI222_X2 i_6_1_882 (.ZN (n_6_1_464), .A1 (n_6_1197), .A2 (slo___n23466), .B1 (n_6_1165)
    , .B2 (slo___n23364), .C1 (slo___n19058), .C2 (n_6_1_483));
INV_X2 i_6_1_881 (.ZN (n_6_2337), .A (n_6_1_464));
BUF_X32 drc_ipo_c29981 (.Z (drc_ipo_n26606), .A (Multiplier[11]));
INV_X2 i_6_1_879 (.ZN (n_6_2336), .A (slo__sro_n16936));
AOI222_X2 slo__sro_c19115 (.ZN (slo__sro_n16920), .A1 (n_6_1261), .A2 (slo___n23274)
    , .B1 (n_6_1229), .B2 (slo___n23359), .C1 (n_6_2338), .C2 (n_6_1_448));
INV_X2 i_6_1_877 (.ZN (n_6_2335), .A (slo__sro_n16886));
NAND2_X1 slo__sro_c7656 (.ZN (slo__sro_n7189), .A1 (n_6_2452), .A2 (n_6_1_588));
INV_X1 i_6_1_875 (.ZN (n_6_2334), .A (CLOCK_slo__sro_n50522));
AOI222_X2 slo__sro_c12404 (.ZN (n_6_1_923), .A1 (n_6_369), .A2 (n_6_1_940), .B1 (n_6_337)
    , .B2 (n_6_1_939), .C1 (n_6_2776), .C2 (CLOCK_sgo__n46937));
INV_X2 i_6_1_873 (.ZN (n_6_2333), .A (slo__sro_n11383));
NAND2_X1 slo__sro_c6400 (.ZN (slo__sro_n6039), .A1 (slo__sro_n6040), .A2 (slo__sro_n6041));
INV_X1 i_6_1_871 (.ZN (slo___n17155), .A (CLOCK_slo__sro_n49772));
NAND2_X1 CLOCK_slo__sro_c66053 (.ZN (CLOCK_slo__sro_n59534), .A1 (CLOCK_sgo__n48020), .A2 (n_6_1777));
BUF_X32 drc_ipo_c29976 (.Z (drc_ipo_n26599), .A (slo__n11938));
AOI222_X2 i_6_1_868 (.ZN (n_6_1_457), .A1 (n_6_1190), .A2 (slo___n23466), .B1 (n_6_1158)
    , .B2 (slo___n23364), .C1 (n_6_2362), .C2 (n_6_1_483));
INV_X1 i_6_1_867 (.ZN (n_6_2330), .A (n_6_1_457));
INV_X1 slo__c42467 (.ZN (slo__n38401), .A (CLOCK_slo__sro_n62783));
INV_X1 i_6_1_865 (.ZN (n_6_2329), .A (n_6_1_456));
NAND2_X1 slo__sro_c15180 (.ZN (slo__sro_n13740), .A1 (n_6_2497), .A2 (n_6_1_623));
BUF_X32 drc_ipo_c29983 (.Z (drc_ipo_n26609), .A (Multiplier[14]));
AND2_X1 slo__sro_c7960 (.ZN (slo__sro_n7478), .A1 (n_6_2544), .A2 (n_6_1_693));
NAND2_X1 slo__sro_c34069 (.ZN (slo__sro_n30504), .A1 (slo__sro_n30505), .A2 (slo__sro_n30506));
NAND2_X1 slo__sro_c7251 (.ZN (slo__sro_n6828), .A1 (slo__sro_n6829), .A2 (slo__sro_n6830));
INV_X1 i_6_1_859 (.ZN (slo___n16361), .A (slo__sro_n6817));
AOI222_X2 i_6_1_858 (.ZN (n_6_1_452), .A1 (n_6_1153), .A2 (slo___n23364), .B1 (n_6_1185)
    , .B2 (slo___n23466), .C1 (slo__n13570), .C2 (n_6_1_483));
NAND2_X1 CLOCK_sgo__sro_c52081 (.ZN (CLOCK_sgo__sro_n47732), .A1 (CLOCK_sgo__sro_n47733), .A2 (CLOCK_sgo__sro_n47734));
AOI222_X1 i_6_1_856 (.ZN (n_6_1_451), .A1 (n_6_1152), .A2 (slo___n23364), .B1 (n_6_1184)
    , .B2 (slo___n23466), .C1 (n_6_2356), .C2 (n_6_1_483));
INV_X1 i_6_1_855 (.ZN (n_6_2324), .A (n_6_1_451));
NOR2_X4 i_6_1_854 (.ZN (n_6_1_450), .A1 (n_6_1_1135), .A2 (Multiplicand[19]));
NOR2_X1 i_6_1_853 (.ZN (n_6_1_449), .A1 (Multiplicand[20]), .A2 (n_6_1_1134));
NOR2_X4 i_6_1_852 (.ZN (n_6_1_448), .A1 (slo___n23274), .A2 (n_6_1_449));
AND2_X1 i_6_1_851 (.ZN (n_6_1_447), .A1 (n_6_2354), .A2 (n_6_1_448));
AOI221_X2 i_6_1_850 (.ZN (n_6_1_446), .A (n_6_1_447), .B1 (n_6_1246), .B2 (slo___n23359)
    , .C1 (n_6_1278), .C2 (slo___n23274));
INV_X2 i_6_1_849 (.ZN (n_6_2323), .A (n_6_1_446));
AOI221_X2 i_6_1_848 (.ZN (n_6_1_445), .A (n_6_1_447), .B1 (n_6_1245), .B2 (slo___n23359)
    , .C1 (n_6_1277), .C2 (slo___n23274));
INV_X2 i_6_1_847 (.ZN (n_6_2322), .A (n_6_1_445));
AOI221_X2 slo__sro_c30790 (.ZN (slo__sro_n27391), .A (slo__sro_n27392), .B1 (n_6_338)
    , .B2 (n_6_1_939), .C1 (n_6_370), .C2 (n_6_1_940));
INV_X2 slo__c46251 (.ZN (n_6_1_542), .A (slo__n41747));
NAND2_X2 slo__sro_c43099 (.ZN (slo__sro_n38941), .A1 (slo__sro_n38942), .A2 (slo__sro_n38943));
INV_X1 i_6_1_843 (.ZN (n_6_2320), .A (CLOCK_sgo__sro_n47835));
AOI222_X1 slo__sro_c11308 (.ZN (n_6_1_73), .A1 (n_6_1863), .A2 (n_6_1_99), .B1 (n_6_1895)
    , .B2 (n_6_1_100), .C1 (n_6_2022), .C2 (n_6_1_98));
INV_X2 i_6_1_841 (.ZN (n_6_2319), .A (n_6_1_442));
NAND2_X1 slo__sro_c6974 (.ZN (slo__sro_n6579), .A1 (n_6_2111), .A2 (n_6_1_203));
INV_X2 i_6_1_839 (.ZN (n_6_2318), .A (slo__sro_n6503));
AND2_X1 slo__sro_c12931 (.ZN (slo__sro_n11858), .A1 (n_6_2792), .A2 (n_6_1_973));
INV_X2 i_6_1_837 (.ZN (n_6_2317), .A (n_6_1_440));
AOI222_X2 i_6_1_836 (.ZN (n_6_1_439), .A1 (n_6_1271), .A2 (slo___n23274), .B1 (n_6_1239)
    , .B2 (slo___n23359), .C1 (n_6_2348), .C2 (n_6_1_448));
INV_X1 i_6_1_835 (.ZN (n_6_2316), .A (n_6_1_439));
AND2_X1 slo__sro_c5999 (.ZN (slo__sro_n5679), .A1 (n_6_2370), .A2 (n_6_1_483));
INV_X1 i_6_1_833 (.ZN (n_6_2315), .A (n_6_1_438));
NAND2_X1 slo__sro_c6746 (.ZN (slo__sro_n6368), .A1 (n_6_2058), .A2 (n_6_1_133));
INV_X2 i_6_1_831 (.ZN (n_6_2314), .A (CLOCK_slo__sro_n55019));
AOI222_X2 i_6_1_830 (.ZN (n_6_1_436), .A1 (n_6_1268), .A2 (slo___n23274), .B1 (n_6_1236)
    , .B2 (slo___n23359), .C1 (n_6_2345), .C2 (n_6_1_448));
INV_X1 i_6_1_829 (.ZN (n_6_2313), .A (n_6_1_436));
NAND2_X1 CLOCK_slo__sro_c58032 (.ZN (CLOCK_slo__sro_n52915), .A1 (CLOCK_slo__sro_n52916), .A2 (CLOCK_slo__sro_n52917));
INV_X2 i_6_1_827 (.ZN (n_6_2312), .A (CLOCK_slo__sro_n52466));
AOI222_X2 i_6_1_826 (.ZN (n_6_1_434), .A1 (n_6_1266), .A2 (slo___n23274), .B1 (n_6_1234)
    , .B2 (slo___n23359), .C1 (n_6_2343), .C2 (n_6_1_448));
INV_X2 i_6_1_825 (.ZN (n_6_2311), .A (n_6_1_434));
AOI222_X2 i_6_1_824 (.ZN (n_6_1_433), .A1 (n_6_1265), .A2 (slo___n23274), .B1 (n_6_1233)
    , .B2 (slo___n23359), .C1 (n_6_2342), .C2 (n_6_1_448));
INV_X1 i_6_1_823 (.ZN (n_6_2310), .A (n_6_1_433));
NAND2_X1 slo__sro_c4520 (.ZN (slo__sro_n4341), .A1 (n_6_2523), .A2 (n_6_1_658));
INV_X1 i_6_1_821 (.ZN (n_6_2309), .A (slo__sro_n4312));
AOI21_X2 CLOCK_slo__sro_c57129 (.ZN (CLOCK_slo__sro_n52126), .A (n_6_1_482), .B1 (n_6_1181), .B2 (slo___n23364));
INV_X2 i_6_1_819 (.ZN (n_6_2308), .A (slo__sro_n39122));
AND2_X1 slo__sro_c9844 (.ZN (slo__sro_n9165), .A1 (n_6_2560), .A2 (n_6_1_693));
INV_X1 i_6_1_817 (.ZN (n_6_2307), .A (slo__sro_n9138));
AOI222_X2 slo__sro_c19137 (.ZN (slo__sro_n16936), .A1 (n_6_1196), .A2 (slo___n23466)
    , .B1 (n_6_1164), .B2 (slo___n23364), .C1 (n_6_2368), .C2 (n_6_1_483));
INV_X2 i_6_1_815 (.ZN (n_6_2306), .A (slo__sro_n16920));
NAND2_X1 slo__sro_c7323 (.ZN (slo__sro_n6899), .A1 (n_6_2190), .A2 (n_6_1_273));
INV_X2 i_6_1_813 (.ZN (n_6_2305), .A (slo__sro_n6827));
NAND2_X1 CLOCK_slo__sro_c65160 (.ZN (CLOCK_slo__sro_n58709), .A1 (CLOCK_slo__sro_n58710), .A2 (slo__sro_n35145));
INV_X2 i_6_1_811 (.ZN (n_6_2304), .A (slo__sro_n40936));
NAND2_X1 slo__sro_c25320 (.ZN (slo__sro_n22113), .A1 (n_6_2626), .A2 (n_6_1_763));
INV_X1 i_6_1_809 (.ZN (n_6_2303), .A (slo__sro_n19997));
AOI222_X1 slo__sro_c10421 (.ZN (slo__sro_n9701), .A1 (n_6_1224), .A2 (slo___n23359)
    , .B1 (n_6_1256), .B2 (slo___n23274), .C1 (n_6_2333), .C2 (n_6_1_448));
INV_X1 i_6_1_807 (.ZN (n_6_2302), .A (slo__sro_n20285));
NAND2_X1 slo__sro_c10432 (.ZN (slo__sro_n9712), .A1 (n_6_1_975), .A2 (n_6_292));
INV_X1 i_6_1_805 (.ZN (n_6_2301), .A (slo__sro_n9701));
INV_X1 slo__c20154 (.ZN (slo__n17720), .A (slo__sro_n31816));
INV_X1 i_6_1_803 (.ZN (n_6_2300), .A (slo__sro_n17693));
NAND2_X1 slo__sro_c13377 (.ZN (slo__sro_n12257), .A1 (opt_ipo_n44599), .A2 (n_6_1_728));
INV_X2 i_6_1_801 (.ZN (n_6_2299), .A (slo__sro_n19543));
INV_X1 CLOCK_slo__sro_c54582 (.ZN (CLOCK_slo__sro_n49913), .A (n_6_1_237));
INV_X1 i_6_1_799 (.ZN (n_6_2298), .A (slo__sro_n6038));
NAND2_X1 slo__sro_c5535 (.ZN (slo__sro_n5270), .A1 (n_6_2681), .A2 (CLOCK_sgo__n46922));
INV_X1 i_6_1_797 (.ZN (n_6_2297), .A (slo__sro_n16910));
AOI222_X2 i_6_1_796 (.ZN (n_6_1_419), .A1 (n_6_1251), .A2 (slo___n23274), .B1 (n_6_1219)
    , .B2 (slo___n23359), .C1 (CLOCK_opt_ipo_n46265), .C2 (n_6_1_448));
AOI21_X1 CLOCK_sgo__sro_c51535 (.ZN (slo__sro_n28562), .A (CLOCK_sgo__sro_n47286)
    , .B1 (n_6_1385), .B2 (n_6_1_380));
NAND2_X1 slo__sro_c6218 (.ZN (slo__sro_n5878), .A1 (n_6_2148), .A2 (n_6_1_238));
INV_X2 i_6_1_793 (.ZN (n_6_2295), .A (slo__sro_n5865));
INV_X1 slo__c20631 (.ZN (slo__n18084), .A (CLOCK_slo__sro_n49022));
INV_X2 i_6_1_791 (.ZN (n_6_2294), .A (slo__sro_n18042));
NAND2_X1 slo__sro_c25675 (.ZN (slo__sro_n22433), .A1 (opt_ipo_n24503), .A2 (n_6_1_973));
INV_X2 i_6_1_789 (.ZN (n_6_2293), .A (slo__sro_n22415));
NOR2_X4 i_6_1_788 (.ZN (n_6_1_415), .A1 (n_6_1_1136), .A2 (Multiplicand[20]));
NOR2_X1 i_6_1_787 (.ZN (CLOCK_slo__n49140), .A1 (Multiplicand[21]), .A2 (n_6_1_1135));
NOR2_X4 i_6_1_786 (.ZN (n_6_1_413), .A1 (slo___n43257), .A2 (n_6_1_414));
AND2_X1 i_6_1_785 (.ZN (n_6_1_412), .A1 (n_6_2323), .A2 (n_6_1_413));
AOI221_X1 i_6_1_784 (.ZN (n_6_1_411), .A (n_6_1_412), .B1 (n_6_1310), .B2 (n_6_1_414)
    , .C1 (n_6_1342), .C2 (slo___n43257));
INV_X2 i_6_1_783 (.ZN (n_6_2292), .A (n_6_1_411));
INV_X1 CLOCK_slo__sro_c59221 (.ZN (CLOCK_slo__sro_n53931), .A (CLOCK_slo__sro_n53932));
INV_X1 i_6_1_781 (.ZN (n_6_2291), .A (CLOCK_slo__sro_n53892));
AND2_X1 slo__sro_c12686 (.ZN (slo__sro_n11641), .A1 (n_6_2414), .A2 (n_6_1_518));
NAND2_X1 slo__sro_c32239 (.ZN (slo__sro_n28775), .A1 (slo__sro_n28776), .A2 (slo__sro_n28777));
AND2_X1 slo__sro_c11290 (.ZN (slo__sro_n10458), .A1 (n_6_2351), .A2 (n_6_1_448));
INV_X2 i_6_1_777 (.ZN (n_6_2289), .A (slo__sro_n10426));
AOI221_X2 slo__sro_c22694 (.ZN (slo__sro_n19695), .A (slo__sro_n19696), .B1 (n_6_1174)
    , .B2 (slo___n23364), .C1 (n_6_1206), .C2 (slo___n23466));
INV_X2 i_6_1_775 (.ZN (slo___n13086), .A (slo__sro_n19567));
NAND2_X1 slo__sro_c12865 (.ZN (slo__sro_n11799), .A1 (opt_ipo_n24190), .A2 (CLOCK_sgo__n46950));
INV_X2 i_6_1_773 (.ZN (n_6_2287), .A (slo__sro_n11754));
AOI222_X2 slo__sro_c13868 (.ZN (slo__sro_n12647), .A1 (n_6_1743), .A2 (n_6_1_169)
    , .B1 (n_6_1775), .B2 (CLOCK_sgo__n48020), .C1 (n_6_2092), .C2 (n_6_1_168));
INV_X2 i_6_1_771 (.ZN (n_6_2286), .A (slo__sro_n12568));
NAND2_X1 slo__sro_c6454 (.ZN (slo__sro_n6090), .A1 (n_6_2469), .A2 (n_6_1_588));
INV_X1 i_6_1_769 (.ZN (n_6_2285), .A (slo__sro_n20680));
NAND2_X1 slo__sro_c37267 (.ZN (slo__sro_n33598), .A1 (n_6_2132), .A2 (n_6_1_203));
INV_X2 i_6_1_767 (.ZN (n_6_2284), .A (slo__sro_n33373));
AND2_X1 slo__sro_c5273 (.ZN (slo__sro_n5027), .A1 (opt_ipo_n24063), .A2 (n_6_1_378));
INV_X1 i_6_1_765 (.ZN (n_6_2283), .A (CLOCK_slo__sro_n61394));
NAND2_X1 slo__sro_c22419 (.ZN (slo__sro_n19439), .A1 (n_6_1_763), .A2 (n_6_2611));
AOI222_X1 slo__sro_c41976 (.ZN (slo__sro_n37999), .A1 (n_6_1513), .A2 (slo___n23247)
    , .B1 (n_6_1481), .B2 (n_6_1_309), .C1 (n_6_2210), .C2 (n_6_1_308));
INV_X1 slo__sro_c15617 (.ZN (slo__sro_n14084), .A (slo__sro_n4923));
INV_X1 i_6_1_761 (.ZN (n_6_2281), .A (slo__sro_n40459));
NAND2_X1 slo__sro_c34678 (.ZN (slo__sro_n31089), .A1 (n_6_2391), .A2 (n_6_1_518));
INV_X2 i_6_1_759 (.ZN (n_6_2280), .A (slo__sro_n31050));
INV_X2 CLOCK_slo__c59027 (.ZN (CLOCK_slo__n53754), .A (slo__sro_n9753));
INV_X1 i_6_1_757 (.ZN (slo__n32747), .A (n_6_1_398));
AOI222_X1 i_6_1_756 (.ZN (n_6_1_397), .A1 (n_6_1328), .A2 (slo___n43257), .B1 (n_6_1296)
    , .B2 (n_6_1_414), .C1 (n_6_2310), .C2 (n_6_1_413));
INV_X2 i_6_1_755 (.ZN (n_6_2278), .A (n_6_1_397));
AOI21_X2 slo__sro_c41071 (.ZN (n_6_1_756), .A (slo__sro_n37209), .B1 (n_6_697), .B2 (n_6_1_765));
INV_X1 i_6_1_753 (.ZN (n_6_2277), .A (n_6_1_396));
NAND2_X1 slo__sro_c7249 (.ZN (slo__sro_n6830), .A1 (n_6_2337), .A2 (n_6_1_448));
INV_X1 i_6_1_751 (.ZN (spw__n67799), .A (slo__sro_n6790));
AOI222_X2 i_6_1_750 (.ZN (n_6_1_394), .A1 (n_6_1325), .A2 (slo___n43257), .B1 (n_6_1293)
    , .B2 (n_6_1_414), .C1 (slo__n12014), .C2 (n_6_1_413));
INV_X1 i_6_1_749 (.ZN (n_6_2275), .A (n_6_1_394));
NAND2_X1 CLOCK_slo__sro_c65838 (.ZN (CLOCK_slo__sro_n59345), .A1 (n_6_2498), .A2 (n_6_1_623));
INV_X2 i_6_1_747 (.ZN (n_6_2274), .A (CLOCK_slo__sro_n64180));
INV_X1 CLOCK_slo__c67283 (.ZN (n_6_1_74), .A (CLOCK_slo__sro_n64636));
INV_X2 i_6_1_745 (.ZN (n_6_2273), .A (slo__sro_n37974));
AOI222_X1 i_6_1_744 (.ZN (slo__n28539), .A1 (n_6_1322), .A2 (slo___n43257), .B1 (n_6_1290)
    , .B2 (n_6_1_414), .C1 (n_6_2304), .C2 (n_6_1_413));
NAND2_X1 slo__sro_c32013 (.ZN (slo__sro_n28564), .A1 (slo__n28538), .A2 (n_6_1_378));
NAND2_X1 slo__mro_c35227 (.ZN (slo__mro_n31601), .A1 (n_6_1562), .A2 (n_6_1_274));
INV_X1 i_6_1_741 (.ZN (n_6_2271), .A (slo__sro_n31234));
NAND2_X1 slo__sro_c10380 (.ZN (slo__sro_n9673), .A1 (n_6_2795), .A2 (n_6_1_973));
INV_X1 i_6_1_739 (.ZN (n_6_2270), .A (slo__sro_n9559));
NAND2_X1 slo__sro_c6613 (.ZN (slo__sro_n6240), .A1 (slo__sro_n6241), .A2 (slo__sro_n6242));
INV_X1 i_6_1_737 (.ZN (n_6_2269), .A (slo__sro_n6191));
AND2_X2 CLOCK_slo__sro_c66167 (.ZN (CLOCK_slo__sro_n59641), .A1 (n_6_1455), .A2 (n_6_1_345));
INV_X1 i_6_1_735 (.ZN (n_6_2268), .A (slo__sro_n6651));
NAND2_X1 slo__sro_c33190 (.ZN (slo__sro_n29677), .A1 (n_6_2804), .A2 (n_6_1_973));
INV_X4 i_6_1_733 (.ZN (n_6_2267), .A (slo__sro_n29650));
INV_X1 slo__sro_c10032 (.ZN (slo__sro_n9342), .A (slo__sro_n9343));
INV_X2 i_6_1_731 (.ZN (n_6_2266), .A (slo__sro_n9242));
AND2_X1 slo__sro_c7481 (.ZN (slo__sro_n7038), .A1 (n_6_2229), .A2 (n_6_1_308));
CLKBUF_X2 CLOCK_sgo__c52408 (.Z (CLOCK_sgo__n48011), .A (n_6_1_99));
NAND2_X1 slo__sro_c7091 (.ZN (slo__sro_n6691), .A1 (n_6_1_413), .A2 (n_6_2297));
NAND2_X2 CLOCK_sgo__sro_c51437 (.ZN (CLOCK_sgo__sro_n47210), .A1 (CLOCK_sgo__sro_n47211), .A2 (CLOCK_sgo__sro_n47212));
AOI222_X1 CLOCK_slo__sro_c61893 (.ZN (slo__sro_n12465), .A1 (n_6_723), .A2 (n_6_1_729)
    , .B1 (n_6_755), .B2 (n_6_1_730), .C1 (n_6_2592), .C2 (n_6_1_728));
INV_X2 i_6_1_725 (.ZN (n_6_2263), .A (slo__sro_n18343));
AOI222_X2 i_6_1_724 (.ZN (n_6_1_381), .A1 (n_6_1312), .A2 (slo___n43257), .B1 (n_6_1280)
    , .B2 (n_6_1_414), .C1 (n_6_2294), .C2 (n_6_1_413));
INV_X2 i_6_1_723 (.ZN (n_6_2262), .A (n_6_1_381));
NOR2_X1 i_6_1_722 (.ZN (slo__n23398), .A1 (n_6_1_1137), .A2 (Multiplicand[21]));
NOR2_X1 i_6_1_721 (.ZN (slo__n23298), .A1 (Multiplicand[22]), .A2 (n_6_1_1136));
NOR2_X4 i_6_1_720 (.ZN (n_6_1_378), .A1 (n_6_1_380), .A2 (n_6_1_379));
AND2_X1 i_6_1_719 (.ZN (n_6_1_377), .A1 (n_6_2292), .A2 (n_6_1_378));
AOI221_X2 i_6_1_718 (.ZN (n_6_1_376), .A (n_6_1_377), .B1 (n_6_1374), .B2 (n_6_1_379)
    , .C1 (n_6_1406), .C2 (n_6_1_380));
INV_X1 i_6_1_717 (.ZN (n_6_2261), .A (n_6_1_376));
AOI221_X2 i_6_1_716 (.ZN (n_6_1_375), .A (n_6_1_377), .B1 (n_6_1373), .B2 (n_6_1_379)
    , .C1 (n_6_1405), .C2 (n_6_1_380));
INV_X2 i_6_1_715 (.ZN (n_6_2260), .A (n_6_1_375));
AND2_X1 slo__sro_c10696 (.ZN (slo__sro_n9948), .A1 (n_6_2631), .A2 (n_6_1_763));
INV_X2 i_6_1_713 (.ZN (n_6_2259), .A (CLOCK_slo__sro_n52632));
NAND2_X1 slo__sro_c5306 (.ZN (slo__sro_n5059), .A1 (slo__n12843), .A2 (n_6_1_308));
INV_X2 i_6_1_711 (.ZN (n_6_2258), .A (CLOCK_sgo__sro_n47798));
NAND2_X1 slo__sro_c10265 (.ZN (slo__sro_n9561), .A1 (n_6_2302), .A2 (n_6_1_413));
INV_X2 i_6_1_709 (.ZN (n_6_2257), .A (slo__sro_n9533));
NAND2_X2 CLOCK_sgo__sro_c51502 (.ZN (CLOCK_sgo__sro_n47261), .A1 (CLOCK_sgo__sro_n47262), .A2 (CLOCK_sgo__sro_n47263));
INV_X1 i_6_1_707 (.ZN (n_6_2256), .A (n_6_1_371));
NAND2_X1 slo__sro_c11415 (.ZN (slo__sro_n10562), .A1 (n_6_2072), .A2 (n_6_1_133));
INV_X2 i_6_1_705 (.ZN (n_6_2255), .A (slo__sro_n34276));
AOI222_X2 i_6_1_704 (.ZN (n_6_1_369), .A1 (n_6_1399), .A2 (n_6_1_380), .B1 (n_6_1367)
    , .B2 (n_6_1_379), .C1 (n_6_2286), .C2 (n_6_1_378));
INV_X2 i_6_1_703 (.ZN (n_6_2254), .A (n_6_1_369));
AOI222_X2 i_6_1_702 (.ZN (n_6_1_368), .A1 (n_6_1398), .A2 (n_6_1_380), .B1 (n_6_1366)
    , .B2 (n_6_1_379), .C1 (n_6_2285), .C2 (n_6_1_378));
INV_X2 i_6_1_701 (.ZN (n_6_2253), .A (n_6_1_368));
AOI221_X2 CLOCK_slo__sro_c58256 (.ZN (n_6_1_1018), .A (slo__sro_n17254), .B1 (n_6_135)
    , .B2 (n_6_1_1044), .C1 (n_6_167), .C2 (n_6_1_1045));
INV_X2 i_6_1_699 (.ZN (n_6_2252), .A (CLOCK_slo__sro_n50138));
AOI21_X4 CLOCK_slo__sro_c58457 (.ZN (slo__sro_n27726), .A (CLOCK_slo__sro_n53277)
    , .B1 (n_6_1596), .B2 (slo___n23244));
INV_X1 slo__L1_c1_c36128 (.ZN (slo__n32451), .A (slo__sro_n38684));
AOI222_X2 i_6_1_696 (.ZN (n_6_1_365), .A1 (n_6_1395), .A2 (n_6_1_380), .B1 (n_6_1363)
    , .B2 (n_6_1_379), .C1 (opt_ipo_n24727), .C2 (n_6_1_378));
INV_X2 i_6_1_695 (.ZN (n_6_2250), .A (n_6_1_365));
NAND2_X1 slo__sro_c8215 (.ZN (slo__sro_n7708), .A1 (n_6_2587), .A2 (n_6_1_728));
INV_X2 i_6_1_693 (.ZN (n_6_2249), .A (n_6_1_364));
NAND2_X1 slo__sro_c7842 (.ZN (slo__sro_n7371), .A1 (n_6_2483), .A2 (n_6_1_623));
INV_X2 i_6_1_691 (.ZN (n_6_2248), .A (slo__sro_n7306));
AOI222_X1 slo__sro_c14891 (.ZN (spt__n66415), .A1 (n_6_1707), .A2 (slo___n23407), .B1 (n_6_1675)
    , .B2 (slo___n23239), .C1 (n_6_2119), .C2 (n_6_1_203));
INV_X1 i_6_1_689 (.ZN (n_6_2247), .A (slo__sro_n13471));
NAND2_X1 slo__sro_c24827 (.ZN (slo__sro_n21665), .A1 (n_6_2485), .A2 (n_6_1_623));
INV_X1 i_6_1_687 (.ZN (n_6_2246), .A (n_6_1_361));
AND2_X1 slo__sro_c23486 (.ZN (slo__sro_n20420), .A1 (n_6_2531), .A2 (n_6_1_658));
INV_X1 i_6_1_685 (.ZN (n_6_2245), .A (CLOCK_slo__sro_n48812));
AOI222_X2 i_6_1_684 (.ZN (n_6_1_359), .A1 (n_6_1389), .A2 (n_6_1_380), .B1 (n_6_1357)
    , .B2 (n_6_1_379), .C1 (CLOCK_slo___n53904), .C2 (n_6_1_378));
INV_X1 i_6_1_683 (.ZN (n_6_2244), .A (n_6_1_359));
AOI222_X2 i_6_1_682 (.ZN (n_6_1_358), .A1 (n_6_1388), .A2 (n_6_1_380), .B1 (n_6_1356)
    , .B2 (n_6_1_379), .C1 (n_6_2275), .C2 (n_6_1_378));
INV_X2 i_6_1_681 (.ZN (n_6_2243), .A (n_6_1_358));
AOI222_X2 i_6_1_680 (.ZN (n_6_1_357), .A1 (n_6_1387), .A2 (n_6_1_380), .B1 (n_6_1355)
    , .B2 (n_6_1_379), .C1 (n_6_2274), .C2 (n_6_1_378));
INV_X2 i_6_1_679 (.ZN (n_6_2242), .A (n_6_1_357));
NAND2_X1 slo__sro_c4521 (.ZN (slo__sro_n4340), .A1 (n_6_844), .A2 (slo___n23463));
INV_X2 i_6_1_677 (.ZN (n_6_2241), .A (n_6_1_356));
AOI221_X2 slo__sro_c32044 (.ZN (slo__sro_n28591), .A (slo__sro_n28592), .B1 (n_6_910)
    , .B2 (slo___n23367), .C1 (n_6_942), .C2 (n_6_1_625));
INV_X1 i_6_1_675 (.ZN (n_6_2240), .A (slo__sro_n28562));
NAND2_X2 CLOCK_slo__sro_c54306 (.ZN (CLOCK_slo__sro_n49674), .A1 (n_6_1348), .A2 (n_6_1_379));
NAND2_X2 CLOCK_sgo__sro_c52504 (.ZN (CLOCK_sgo__sro_n48086), .A1 (n_6_290), .A2 (n_6_1_975));
NAND2_X1 slo__sro_c23314 (.ZN (slo__sro_n20261), .A1 (n_6_912), .A2 (slo___n23367));
INV_X4 i_6_1_671 (.ZN (n_6_2238), .A (slo__sro_n20146));
NAND2_X1 CLOCK_slo__sro_c54416 (.ZN (CLOCK_slo__sro_n49775), .A1 (n_6_2364), .A2 (n_6_1_483));
INV_X2 i_6_1_669 (.ZN (n_6_2237), .A (CLOCK_slo__sro_n49758));
AOI21_X2 slo__sro_c6315 (.ZN (n_6_1_741), .A (slo__sro_n5963), .B1 (n_6_650), .B2 (n_6_1_764));
INV_X2 i_6_1_667 (.ZN (n_6_2236), .A (slo__sro_n5945));
AOI221_X2 slo__sro_c10121 (.ZN (slo__n27411), .A (slo__sro_n9421), .B1 (n_6_1881)
    , .B2 (CLOCK_sgo__n48011), .C1 (n_6_1913), .C2 (n_6_1_100));
INV_X1 i_6_1_665 (.ZN (n_6_2235), .A (CLOCK_slo__sro_n49672));
AOI21_X1 CLOCK_slo__sro_c57684 (.ZN (CLOCK_slo__sro_n52592), .A (CLOCK_slo__sro_n52593)
    , .B1 (n_6_1613), .B2 (slo___n23215));
INV_X2 i_6_1_663 (.ZN (n_6_2234), .A (n_6_1_349));
NAND2_X1 slo__sro_c10031 (.ZN (slo__sro_n9343), .A1 (n_6_2769), .A2 (CLOCK_sgo__n46937));
INV_X2 i_6_1_661 (.ZN (n_6_2233), .A (slo__sro_n36308));
AOI222_X1 i_6_1_660 (.ZN (n_6_1_347), .A1 (n_6_1377), .A2 (n_6_1_380), .B1 (n_6_1345)
    , .B2 (n_6_1_379), .C1 (CLOCK_opt_ipo_n45803), .C2 (n_6_1_378));
INV_X1 i_6_1_659 (.ZN (n_6_2232), .A (n_6_1_347));
AOI222_X1 i_6_1_658 (.ZN (n_6_1_346), .A1 (n_6_1376), .A2 (n_6_1_380), .B1 (n_6_1344)
    , .B2 (n_6_1_379), .C1 (n_6_2263), .C2 (n_6_1_378));
INV_X1 i_6_1_657 (.ZN (n_6_2231), .A (n_6_1_346));
NOR2_X1 i_6_1_656 (.ZN (slo__n23445), .A1 (n_6_1_1138), .A2 (Multiplicand[22]));
NOR2_X4 i_6_1_655 (.ZN (n_6_1_344), .A1 (Multiplicand[23]), .A2 (n_6_1_1137));
NOR2_X4 i_6_1_654 (.ZN (n_6_1_343), .A1 (n_6_1_345), .A2 (slo___n23229));
AND2_X1 i_6_1_653 (.ZN (n_6_1_342), .A1 (n_6_2261), .A2 (n_6_1_343));
AOI221_X2 i_6_1_652 (.ZN (n_6_1_341), .A (n_6_1_342), .B1 (n_6_1438), .B2 (slo___n23229)
    , .C1 (n_6_1470), .C2 (n_6_1_345));
INV_X2 i_6_1_651 (.ZN (n_6_2230), .A (n_6_1_341));
AOI221_X2 i_6_1_650 (.ZN (n_6_1_340), .A (n_6_1_342), .B1 (n_6_1437), .B2 (slo___n23229)
    , .C1 (n_6_1469), .C2 (n_6_1_345));
INV_X2 i_6_1_649 (.ZN (n_6_2229), .A (n_6_1_340));
AOI221_X1 slo__sro_c10553 (.ZN (n_6_1_549), .A (slo__sro_n9815), .B1 (n_6_1052), .B2 (n_6_1_554)
    , .C1 (n_6_1084), .C2 (slo___n23457));
INV_X2 i_6_1_647 (.ZN (n_6_2228), .A (CLOCK_slo__mro_n51371));
NAND2_X1 slo__sro_c34641 (.ZN (slo__sro_n31053), .A1 (n_6_2312), .A2 (n_6_1_413));
INV_X1 i_6_1_645 (.ZN (slo___n15724), .A (slo__sro_n19751));
NAND2_X1 slo__sro_c3093 (.ZN (slo__sro_n3059), .A1 (n_6_2185), .A2 (n_6_1_273));
AOI21_X2 slo__c17659 (.ZN (slo__n15804), .A (slo__sro_n4845), .B1 (n_6_1653), .B2 (drc_ipo_n26601));
INV_X4 i_6_1_641 (.ZN (n_6_2225), .A (slo__sro_n21436));
AND2_X1 CLOCK_slo__sro_c65956 (.ZN (CLOCK_slo__sro_n59448), .A1 (n_6_2223), .A2 (n_6_1_308));
INV_X2 i_6_1_639 (.ZN (n_6_2224), .A (n_6_1_335));
AND2_X1 slo__sro_c10552 (.ZN (slo__sro_n9815), .A1 (n_6_2446), .A2 (n_6_1_553));
INV_X1 i_6_1_637 (.ZN (n_6_2223), .A (slo__sro_n9753));
NAND2_X1 slo__sro_c9925 (.ZN (slo__sro_n9245), .A1 (n_6_1_413), .A2 (n_6_2298));
INV_X2 i_6_1_635 (.ZN (n_6_2222), .A (slo__sro_n9194));
AND2_X1 slo__sro_c22693 (.ZN (slo__sro_n19696), .A1 (n_6_2378), .A2 (n_6_1_483));
INV_X4 i_6_1_633 (.ZN (n_6_2221), .A (slo__sro_n19673));
BUF_X32 slo__c5176 (.Z (slo__n4932), .A (n_6_7));
INV_X2 i_6_1_631 (.ZN (n_6_2220), .A (slo__sro_n14081));
INV_X1 CLOCK_slo__sro_c54227 (.ZN (CLOCK_slo__sro_n49605), .A (slo__sro_n8742));
INV_X1 i_6_1_629 (.ZN (n_6_2219), .A (n_6_1_330));
NAND2_X1 slo__sro_c38938 (.ZN (slo__sro_n35272), .A1 (n_6_1_1045), .A2 (n_6_164));
AOI21_X4 slo__sro_c41787 (.ZN (n_6_1_894), .A (slo__sro_n37841), .B1 (n_6_407), .B2 (n_6_1_904));
AOI222_X2 i_6_1_626 (.ZN (n_6_1_328), .A1 (n_6_1457), .A2 (n_6_1_345), .B1 (n_6_1425)
    , .B2 (slo___n23229), .C1 (n_6_2249), .C2 (n_6_1_343));
INV_X1 i_6_1_625 (.ZN (n_6_2217), .A (n_6_1_328));
INV_X2 slo__c40377 (.ZN (slo__n36610), .A (slo__sro_n5678));
INV_X2 i_6_1_623 (.ZN (n_6_2216), .A (slo__sro_n36088));
NAND2_X1 slo__sro_c7291 (.ZN (slo__sro_n6872), .A1 (n_6_2376), .A2 (n_6_1_483));
INV_X2 i_6_1_621 (.ZN (n_6_2215), .A (slo__sro_n6762));
AOI222_X2 i_6_1_620 (.ZN (n_6_1_325), .A1 (n_6_1454), .A2 (n_6_1_345), .B1 (n_6_1422)
    , .B2 (slo___n23229), .C1 (n_6_2246), .C2 (n_6_1_343));
INV_X2 i_6_1_619 (.ZN (n_6_2214), .A (n_6_1_325));
AOI222_X2 i_6_1_618 (.ZN (n_6_1_324), .A1 (n_6_1453), .A2 (n_6_1_345), .B1 (n_6_1421)
    , .B2 (slo___n23229), .C1 (n_6_2245), .C2 (n_6_1_343));
INV_X1 i_6_1_617 (.ZN (n_6_2213), .A (n_6_1_324));
AOI221_X2 slo__sro_c4040 (.ZN (slo__sro_n3904), .A (slo__sro_n3905), .B1 (n_6_1495)
    , .B2 (n_6_1_309), .C1 (n_6_1527), .C2 (slo___n23247));
INV_X2 i_6_1_615 (.ZN (n_6_2212), .A (slo__sro_n3860));
NAND2_X1 CLOCK_slo__sro_c54786 (.ZN (CLOCK_slo__sro_n50098), .A1 (n_6_1450), .A2 (n_6_1_345));
INV_X2 i_6_1_613 (.ZN (n_6_2211), .A (CLOCK_slo__sro_n50082));
NAND2_X1 slo__sro_c5369 (.ZN (slo__sro_n5120), .A1 (n_6_1_763), .A2 (n_6_2622));
INV_X2 i_6_1_611 (.ZN (n_6_2210), .A (CLOCK_slo__sro_n50096));
AOI222_X2 i_6_1_610 (.ZN (n_6_1_320), .A1 (n_6_1449), .A2 (n_6_1_345), .B1 (n_6_1417)
    , .B2 (slo___n23229), .C1 (n_6_2241), .C2 (n_6_1_343));
INV_X2 i_6_1_609 (.ZN (n_6_2209), .A (n_6_1_320));
INV_X1 slo__sro_c26503 (.ZN (slo__sro_n23159), .A (slo__sro_n23160));
INV_X4 i_6_1_607 (.ZN (n_6_2208), .A (CLOCK_slo__sro_n53257));
INV_X1 slo__sro_c13472 (.ZN (slo__sro_n12328), .A (slo__sro_n12329));
INV_X4 i_6_1_605 (.ZN (n_6_2207), .A (slo__sro_n12224));
NOR2_X1 slo__sro_c44283 (.ZN (slo__sro_n39888), .A1 (slo__sro_n8356), .A2 (slo__sro_n39889));
INV_X1 i_6_1_603 (.ZN (n_6_2206), .A (slo__sro_n39597));
AOI21_X2 slo__sro_c7052 (.ZN (slo__sro_n6651), .A (slo__sro_n6652), .B1 (n_6_1318), .B2 (slo___n43257));
INV_X2 i_6_1_601 (.ZN (n_6_2205), .A (slo__sro_n40007));
NAND2_X1 slo__sro_c25840 (.ZN (slo__sro_n22580), .A1 (n_6_2113), .A2 (n_6_1_203));
INV_X2 i_6_1_599 (.ZN (n_6_2204), .A (CLOCK_slo__sro_n55084));
AOI222_X2 i_6_1_598 (.ZN (n_6_1_314), .A1 (n_6_1443), .A2 (n_6_1_345), .B1 (n_6_1411)
    , .B2 (slo___n23229), .C1 (n_6_2235), .C2 (n_6_1_343));
INV_X2 i_6_1_597 (.ZN (n_6_2203), .A (n_6_1_314));
NAND2_X1 slo__sro_c42875 (.ZN (slo__sro_n38746), .A1 (n_6_848), .A2 (slo___n23463));
INV_X2 i_6_1_595 (.ZN (n_6_2202), .A (slo__sro_n38408));
NAND2_X1 slo__sro_c7075 (.ZN (slo__sro_n6676), .A1 (n_6_1_413), .A2 (CLOCK_opt_ipo_n45807));
NAND2_X1 CLOCK_slo__sro_c68124 (.ZN (CLOCK_slo__sro_n61349), .A1 (n_6_2853), .A2 (CLOCK_sgo__n46945));
AOI222_X1 i_6_1_592 (.ZN (n_6_1_311), .A1 (n_6_1440), .A2 (n_6_1_345), .B1 (n_6_1408)
    , .B2 (slo___n23229), .C1 (n_6_2232), .C2 (n_6_1_343));
INV_X1 i_6_1_591 (.ZN (n_6_2200), .A (n_6_1_311));
NOR2_X4 i_6_1_590 (.ZN (n_6_1_310), .A1 (n_6_1_1139), .A2 (Multiplicand[23]));
NOR2_X1 i_6_1_589 (.ZN (slo__n23262), .A1 (Multiplicand[24]), .A2 (n_6_1_1138));
NOR2_X4 i_6_1_588 (.ZN (n_6_1_308), .A1 (slo___n23247), .A2 (n_6_1_309));
AND2_X1 i_6_1_587 (.ZN (n_6_1_307), .A1 (n_6_2230), .A2 (n_6_1_308));
AOI221_X2 i_6_1_586 (.ZN (n_6_1_306), .A (n_6_1_307), .B1 (n_6_1502), .B2 (n_6_1_309)
    , .C1 (n_6_1534), .C2 (slo___n23247));
INV_X2 i_6_1_585 (.ZN (n_6_2199), .A (n_6_1_306));
AOI221_X2 i_6_1_584 (.ZN (spt__n66340), .A (n_6_1_307), .B1 (n_6_1501), .B2 (n_6_1_309)
    , .C1 (n_6_1533), .C2 (slo___n23247));
INV_X2 i_6_1_583 (.ZN (n_6_2198), .A (n_6_1_305));
AND2_X1 slo__sro_c7554 (.ZN (slo__sro_n7098), .A1 (n_6_2221), .A2 (n_6_1_308));
INV_X1 i_6_1_581 (.ZN (n_6_2197), .A (slo__sro_n7037));
NAND2_X1 slo__sro_c11527 (.ZN (slo__sro_n10652), .A1 (n_6_2073), .A2 (n_6_1_133));
INV_X2 i_6_1_579 (.ZN (n_6_2196), .A (slo__sro_n28283));
AOI21_X2 CLOCK_slo__sro_c53350 (.ZN (CLOCK_slo__sro_n48812), .A (CLOCK_slo__sro_n48813)
    , .B1 (n_6_1390), .B2 (n_6_1_380));
INV_X2 i_6_1_577 (.ZN (n_6_2195), .A (CLOCK_slo__sro_n48784));
NAND2_X1 slo__sro_c17498 (.ZN (slo__sro_n15671), .A1 (opt_ipo_n45121), .A2 (n_6_1_273));
AOI21_X4 CLOCK_sgo__sro_c51366 (.ZN (n_6_1_699), .A (CLOCK_sgo__sro_n47148), .B1 (n_6_707), .B2 (n_6_1_729));
AND2_X1 slo__sro_c22782 (.ZN (slo__sro_n19776), .A1 (slo__sro_n8179), .A2 (n_6_1_553));
INV_X1 i_6_1_573 (.ZN (n_6_2193), .A (slo__sro_n19627));
AND2_X1 slo__sro_c4343 (.ZN (slo__sro_n4176), .A1 (n_6_1_798), .A2 (n_6_2660));
INV_X2 i_6_1_571 (.ZN (n_6_2192), .A (slo__sro_n3904));
NAND2_X1 slo__sro_c6529 (.ZN (slo__sro_n6163), .A1 (n_6_1_308), .A2 (n_6_2207));
INV_X2 i_6_1_569 (.ZN (n_6_2191), .A (CLOCK_slo__sro_n59447));
NAND2_X2 slo__sro_c14705 (.ZN (slo__sro_n13356), .A1 (n_6_1751), .A2 (n_6_1_169));
INV_X2 i_6_1_567 (.ZN (n_6_2190), .A (slo__sro_n13332));
CLKBUF_X1 slo___L1_c1_c7582 (.Z (n_6_2388), .A (CLOCK_opt_ipo_n45825));
INV_X2 i_6_1_565 (.ZN (n_6_2189), .A (CLOCK_slo__sro_n51060));
NAND2_X1 slo__sro_c32238 (.ZN (slo__sro_n28776), .A1 (n_6_1_765), .A2 (n_6_692));
INV_X1 i_6_1_563 (.ZN (slo___n17633), .A (n_6_1_295));
AOI222_X2 i_6_1_562 (.ZN (n_6_1_294), .A1 (n_6_1522), .A2 (slo___n23247), .B1 (n_6_1490)
    , .B2 (n_6_1_309), .C1 (slo__n39406), .C2 (n_6_1_308));
INV_X1 i_6_1_561 (.ZN (n_6_2187), .A (n_6_1_294));
AOI222_X2 i_6_1_560 (.ZN (n_6_1_293), .A1 (n_6_1521), .A2 (slo___n23247), .B1 (n_6_1489)
    , .B2 (n_6_1_309), .C1 (opt_ipo_n24721), .C2 (n_6_1_308));
INV_X2 i_6_1_559 (.ZN (n_6_2186), .A (n_6_1_293));
INV_X1 CLOCK_slo__sro_c55007 (.ZN (CLOCK_slo__sro_n50303), .A (slo__sro_n12506));
INV_X2 i_6_1_557 (.ZN (n_6_2185), .A (CLOCK_slo__sro_n50224));
INV_X2 slo__c14054 (.ZN (slo__n12811), .A (slo__sro_n7515));
INV_X2 i_6_1_555 (.ZN (n_6_2184), .A (slo__sro_n12743));
NAND2_X1 slo__sro_c22564 (.ZN (slo__sro_n19569), .A1 (n_6_1306), .A2 (n_6_1_414));
INV_X1 i_6_1_553 (.ZN (n_6_2183), .A (slo__sro_n29380));
AND2_X1 slo__sro_c5324 (.ZN (slo__sro_n5075), .A1 (n_6_2242), .A2 (n_6_1_343));
INV_X2 i_6_1_551 (.ZN (n_6_2182), .A (slo__sro_n5056));
NAND2_X1 slo__sro_c11255 (.ZN (slo__sro_n10429), .A1 (n_6_1_413), .A2 (opt_ipo_n45132));
INV_X2 i_6_1_549 (.ZN (n_6_2181), .A (n_6_1_288));
AOI21_X2 slo__sro_c14843 (.ZN (slo__sro_n13471), .A (slo__sro_n13472), .B1 (n_6_1392), .B2 (n_6_1_380));
INV_X2 i_6_1_547 (.ZN (n_6_2180), .A (slo__sro_n13461));
AOI222_X2 i_6_1_546 (.ZN (n_6_1_286), .A1 (n_6_1514), .A2 (slo___n23247), .B1 (n_6_1482)
    , .B2 (n_6_1_309), .C1 (n_6_2211), .C2 (n_6_1_308));
INV_X2 i_6_1_545 (.ZN (n_6_2179), .A (n_6_1_286));
NAND2_X1 slo__sro_c42475 (.ZN (slo__sro_n38410), .A1 (slo___n23229), .A2 (n_6_1410));
INV_X1 i_6_1_543 (.ZN (n_6_2178), .A (slo__sro_n37999));
NAND2_X1 slo__sro_c32862 (.ZN (slo__sro_n29363), .A1 (slo__sro_n29364), .A2 (slo__sro_n29365));
INV_X1 i_6_1_541 (.ZN (n_6_2177), .A (slo__sro_n29225));
AOI222_X2 slo__sro_c14302 (.ZN (slo__sro_n13019), .A1 (n_6_1945), .A2 (n_6_1_64), .B1 (n_6_1977)
    , .B2 (n_6_1_65), .C1 (n_6_2009), .C2 (n_6_1_63));
INV_X4 i_6_1_539 (.ZN (n_6_2176), .A (CLOCK_slo__sro_n51885));
AOI222_X2 slo__sro_c6601 (.ZN (slo__sro_n6229), .A1 (n_6_553), .A2 (n_6_1_835), .B1 (n_6_521)
    , .B2 (n_6_1_834), .C1 (n_6_2675), .C2 (CLOCK_sgo__n46922));
NAND2_X1 CLOCK_sgo__sro_c52215 (.ZN (CLOCK_sgo__sro_n47847), .A1 (n_6_1466), .A2 (n_6_1_345));
CLKBUF_X2 CLOCK_sgo__c52417 (.Z (CLOCK_sgo__n48020), .A (n_6_1_170));
INV_X2 i_6_1_535 (.ZN (n_6_2174), .A (n_6_1_281));
NAND2_X1 CLOCK_slo__sro_c59372 (.ZN (CLOCK_slo__sro_n54054), .A1 (n_6_1040), .A2 (n_6_1_554));
INV_X2 i_6_1_533 (.ZN (n_6_2173), .A (n_6_1_280));
NAND2_X1 slo__sro_c23342 (.ZN (slo__sro_n20287), .A1 (n_6_1257), .A2 (slo___n23274));
AOI221_X2 CLOCK_slo__sro_c68066 (.ZN (CLOCK_slo__sro_n61295), .A (CLOCK_slo__sro_n61296)
    , .B1 (n_6_64), .B2 (n_6_1_1079), .C1 (n_6_96), .C2 (n_6_1_1080));
AOI21_X2 slo__sro_c23582 (.ZN (slo__sro_n20506), .A (slo__mro_n33237), .B1 (n_6_1715), .B2 (slo___n23407));
INV_X2 i_6_1_529 (.ZN (n_6_2171), .A (slo__sro_n20472));
AOI21_X2 slo__sro_c40225 (.ZN (slo__sro_n36476), .A (slo__sro_n36477), .B1 (n_6_1064), .B2 (slo___n23457));
INV_X1 i_6_1_527 (.ZN (n_6_2170), .A (slo__sro_n36260));
AOI222_X2 i_6_1_526 (.ZN (n_6_1_276), .A1 (n_6_1504), .A2 (slo___n23247), .B1 (n_6_1472)
    , .B2 (n_6_1_309), .C1 (CLOCK_opt_ipo_n45893), .C2 (n_6_1_308));
INV_X1 i_6_1_525 (.ZN (n_6_2169), .A (n_6_1_276));
NOR2_X4 i_6_1_524 (.ZN (n_6_1_275), .A1 (n_6_1_1140), .A2 (Multiplicand[24]));
NOR2_X1 i_6_1_523 (.ZN (CLOCK_slo__n50420), .A1 (Multiplicand[25]), .A2 (n_6_1_1139));
NOR2_X4 i_6_1_522 (.ZN (n_6_1_273), .A1 (slo___n23244), .A2 (n_6_1_274));
AND2_X1 i_6_1_521 (.ZN (n_6_1_272), .A1 (n_6_2199), .A2 (n_6_1_273));
NAND2_X1 CLOCK_slo__sro_c64709 (.ZN (CLOCK_slo__sro_n58343), .A1 (n_6_1_973), .A2 (opt_ipo_n25120));
INV_X2 i_6_1_519 (.ZN (n_6_2168), .A (CLOCK_slo__sro_n57699));
AOI221_X2 i_6_1_518 (.ZN (n_6_1_270), .A (n_6_1_272), .B1 (n_6_1565), .B2 (n_6_1_274)
    , .C1 (n_6_1597), .C2 (slo___n23244));
INV_X2 i_6_1_517 (.ZN (n_6_2167), .A (n_6_1_270));
INV_X1 slo__sro_c31252 (.ZN (slo__sro_n27837), .A (slo__sro_n27838));
INV_X1 i_6_1_515 (.ZN (n_6_2166), .A (slo__sro_n27726));
AOI222_X2 i_6_1_514 (.ZN (n_6_1_268), .A1 (n_6_1595), .A2 (slo___n23244), .B1 (n_6_1563)
    , .B2 (n_6_1_274), .C1 (n_6_2197), .C2 (n_6_1_273));
INV_X1 i_6_1_513 (.ZN (n_6_2165), .A (n_6_1_268));
NAND2_X1 slo__sro_c7883 (.ZN (slo__sro_n7406), .A1 (slo__sro_n7407), .A2 (slo__sro_n7408));
INV_X2 i_6_1_511 (.ZN (n_6_2164), .A (n_6_1_267));
INV_X1 slo__sro_c38260 (.ZN (slo__sro_n34622), .A (n_6_1_693));
INV_X2 i_6_1_509 (.ZN (n_6_2163), .A (slo__sro_n34553));
NAND2_X1 slo__sro_c17514 (.ZN (slo__sro_n15687), .A1 (CLOCK_slo__n57308), .A2 (n_6_1_273));
INV_X2 i_6_1_507 (.ZN (n_6_2162), .A (slo__sro_n15668));
NAND2_X1 slo__sro_c17530 (.ZN (slo__sro_n15703), .A1 (n_6_2179), .A2 (n_6_1_273));
INV_X4 i_6_1_505 (.ZN (n_6_2161), .A (slo__sro_n15684));
AOI222_X2 slo__sro_c37430 (.ZN (slo__sro_n33755), .A1 (n_6_197), .A2 (n_6_1_1009)
    , .B1 (n_6_229), .B2 (n_6_1_1010), .C1 (n_6_2826), .C2 (CLOCK_sgo__n46950));
INV_X2 i_6_1_503 (.ZN (n_6_2160), .A (slo__sro_n33526));
INV_X1 slo__sro_c16918 (.ZN (slo__sro_n15199), .A (slo__sro_n15200));
INV_X2 i_6_1_501 (.ZN (n_6_2159), .A (CLOCK_slo__sro_n50730));
NAND2_X1 CLOCK_slo__sro_c55856 (.ZN (CLOCK_slo__sro_n51062), .A1 (n_6_1524), .A2 (slo___n23247));
INV_X1 i_6_1_499 (.ZN (n_6_2158), .A (slo__sro_n6897));
NAND2_X2 slo__sro_c24583 (.ZN (slo__sro_n21437), .A1 (slo__sro_n21438), .A2 (slo__sro_n21439));
INV_X4 i_6_1_497 (.ZN (n_6_2157), .A (n_6_1_260));
NAND2_X1 CLOCK_sgo__sro_c51633 (.ZN (CLOCK_sgo__sro_n47371), .A1 (n_6_2141), .A2 (n_6_1_238));
INV_X2 i_6_1_495 (.ZN (slo___n13169), .A (n_6_1_259));
INV_X1 CLOCK_sgo__sro_c51982 (.ZN (CLOCK_sgo__sro_n47665), .A (slo__sro_n10713));
INV_X2 i_6_1_493 (.ZN (n_6_2155), .A (CLOCK_sgo__sro_n47592));
AOI222_X2 i_6_1_492 (.ZN (n_6_1_257), .A1 (n_6_1584), .A2 (slo___n23244), .B1 (n_6_1552)
    , .B2 (n_6_1_274), .C1 (n_6_2186), .C2 (n_6_1_273));
INV_X2 i_6_1_491 (.ZN (n_6_2154), .A (n_6_1_257));
NAND2_X1 slo__sro_c3870 (.ZN (slo__sro_n3751), .A1 (slo__n38240), .A2 (n_6_1_273));
INV_X4 i_6_1_489 (.ZN (n_6_2153), .A (slo__sro_n3056));
INV_X2 slo__c14214 (.ZN (slo__n12943), .A (n_6_1_294));
INV_X1 i_6_1_487 (.ZN (n_6_2152), .A (slo__sro_n12923));
CLKBUF_X1 CLOCK_spw__L1_c1_c73368 (.Z (opt_ipo_n45480), .A (CLOCK_spw__n65836));
INV_X1 i_6_1_485 (.ZN (n_6_2151), .A (slo__sro_n3748));
AOI21_X2 slo__sro_c42477 (.ZN (slo__sro_n38408), .A (slo__sro_n38409), .B1 (n_6_1442), .B2 (n_6_1_345));
BUF_X1 spt__c74536 (.Z (n_6_1_801), .A (spt__n66327));
INV_X2 i_6_1_481 (.ZN (n_6_2149), .A (n_6_1_252));
NAND2_X1 slo__sro_c13761 (.ZN (slo__sro_n12558), .A1 (n_6_2694), .A2 (CLOCK_sgo__n46922));
INV_X2 i_6_1_479 (.ZN (n_6_2148), .A (slo__sro_n12534));
NAND2_X1 slo__sro_c17692 (.ZN (slo__sro_n15831), .A1 (n_6_1742), .A2 (n_6_1_169));
INV_X1 i_6_1_477 (.ZN (n_6_2147), .A (slo__sro_n15700));
AOI21_X2 slo__sro_c21942 (.ZN (slo__sro_n19076), .A (slo__sro_n19077), .B1 (n_6_627), .B2 (n_6_1_800));
INV_X2 i_6_1_475 (.ZN (n_6_2146), .A (slo__sro_n19024));
AOI222_X2 i_6_1_474 (.ZN (n_6_1_248), .A1 (n_6_1575), .A2 (slo___n23244), .B1 (n_6_1543)
    , .B2 (n_6_1_274), .C1 (n_6_2177), .C2 (n_6_1_273));
INV_X2 i_6_1_473 (.ZN (n_6_2145), .A (n_6_1_248));
NAND2_X1 slo__sro_c23378 (.ZN (slo__sro_n20324), .A1 (slo__n35114), .A2 (n_6_1_518));
INV_X1 i_6_1_471 (.ZN (n_6_2144), .A (slo__sro_n32316));
INV_X1 slo__c21475 (.ZN (slo__n18737), .A (slo__sro_n9341));
INV_X2 i_6_1_469 (.ZN (n_6_2143), .A (CLOCK_slo__sro_n57685));
INV_X1 slo__c20879 (.ZN (slo__n18277), .A (slo__sro_n11034));
INV_X2 i_6_1_467 (.ZN (n_6_2142), .A (n_6_1_245));
AOI222_X2 i_6_1_466 (.ZN (n_6_1_244), .A1 (n_6_1571), .A2 (slo___n23244), .B1 (n_6_1539)
    , .B2 (n_6_1_274), .C1 (n_6_2173), .C2 (n_6_1_273));
INV_X2 i_6_1_465 (.ZN (n_6_2141), .A (n_6_1_244));
AND2_X1 CLOCK_sgo__sro_c52037 (.ZN (CLOCK_sgo__sro_n47701), .A1 (n_6_2145), .A2 (n_6_1_238));
INV_X2 i_6_1_463 (.ZN (n_6_2140), .A (n_6_1_243));
AOI222_X2 i_6_1_462 (.ZN (n_6_1_242), .A1 (n_6_1569), .A2 (slo___n23244), .B1 (n_6_1537)
    , .B2 (n_6_1_274), .C1 (n_6_2171), .C2 (n_6_1_273));
INV_X2 i_6_1_461 (.ZN (n_6_2139), .A (n_6_1_242));
AOI222_X1 i_6_1_460 (.ZN (n_6_1_241), .A1 (n_6_1568), .A2 (slo___n23244), .B1 (n_6_1536)
    , .B2 (n_6_1_274), .C1 (n_6_2170), .C2 (n_6_1_273));
INV_X1 i_6_1_459 (.ZN (n_6_2138), .A (n_6_1_241));
NOR2_X4 i_6_1_458 (.ZN (n_6_1_240), .A1 (n_6_1_1141), .A2 (Multiplicand[25]));
NOR2_X4 i_6_1_457 (.ZN (n_6_1_239), .A1 (Multiplicand[26]), .A2 (n_6_1_1140));
NOR2_X4 i_6_1_456 (.ZN (n_6_1_238), .A1 (drc_ipo_n26601), .A2 (slo___n23215));
AND2_X1 i_6_1_455 (.ZN (n_6_1_237), .A1 (n_6_2168), .A2 (n_6_1_238));
NAND2_X1 CLOCK_slo__sro_c54402 (.ZN (CLOCK_slo__sro_n49761), .A1 (n_6_2269), .A2 (n_6_1_378));
INV_X1 i_6_1_453 (.ZN (n_6_2137), .A (n_6_1_236));
INV_X1 CLOCK_slo__sro_c54615 (.ZN (CLOCK_slo__sro_n49939), .A (n_6_2037));
INV_X2 i_6_1_451 (.ZN (n_6_2136), .A (n_6_1_235));
INV_X1 slo__sro_c23759 (.ZN (slo__sro_n20683), .A (slo__sro_n6021));
INV_X4 i_6_1_449 (.ZN (n_6_2135), .A (slo__sro_n32163));
NAND2_X1 slo__sro_c4889 (.ZN (slo__sro_n4673), .A1 (n_6_1_1045), .A2 (n_6_169));
INV_X1 i_6_1_447 (.ZN (n_6_2134), .A (n_6_1_233));
AOI221_X2 slo__sro_c38807 (.ZN (n_6_1_440), .A (slo__sro_n11844), .B1 (n_6_1272), .B2 (slo___n23274)
    , .C1 (n_6_1240), .C2 (slo___n23359));
INV_X2 i_6_1_445 (.ZN (n_6_2133), .A (CLOCK_slo__sro_n58708));
INV_X1 slo__sro_c23914 (.ZN (slo__sro_n20819), .A (n_6_1_798));
INV_X2 i_6_1_443 (.ZN (n_6_2132), .A (n_6_1_231));
AOI221_X2 slo__sro_c5007 (.ZN (slo__sro_n4774), .A (slo__sro_n4775), .B1 (n_6_1110)
    , .B2 (slo___n23277), .C1 (n_6_1142), .C2 (n_6_1_520));
INV_X2 i_6_1_441 (.ZN (slo__n30795), .A (CLOCK_slo__sro_n54099));
AOI21_X1 slo__sro_c14682 (.ZN (slo__sro_n13332), .A (slo__sro_n13333), .B1 (n_6_1525), .B2 (slo___n23247));
INV_X2 i_6_1_439 (.ZN (n_6_2130), .A (slo__sro_n22132));
NAND2_X1 slo__sro_c6914 (.ZN (slo__sro_n6522), .A1 (slo__n13799), .A2 (n_6_2905));
NAND2_X2 CLOCK_sgo__sro_c52163 (.ZN (CLOCK_sgo__sro_n47799), .A1 (CLOCK_sgo__sro_n47800), .A2 (CLOCK_sgo__sro_n47801));
NAND2_X1 slo__sro_c5121 (.ZN (slo__sro_n4883), .A1 (n_6_2404), .A2 (n_6_1_518));
INV_X1 i_6_1_435 (.ZN (n_6_2128), .A (slo__sro_n4844));
AOI222_X2 i_6_1_434 (.ZN (n_6_1_226), .A1 (n_6_1652), .A2 (drc_ipo_n26601), .B1 (n_6_1620)
    , .B2 (slo___n23215), .C1 (n_6_2159), .C2 (n_6_1_238));
INV_X2 i_6_1_433 (.ZN (n_6_2127), .A (n_6_1_226));
NAND2_X1 CLOCK_slo__sro_c63884 (.ZN (CLOCK_slo__sro_n57700), .A1 (CLOCK_slo__sro_n57701), .A2 (CLOCK_slo__sro_n57702));
INV_X2 i_6_1_431 (.ZN (n_6_2126), .A (slo__sro_n15342));
NAND2_X1 slo__sro_c32237 (.ZN (slo__sro_n28777), .A1 (n_6_1_763), .A2 (slo___n12846));
INV_X2 i_6_1_429 (.ZN (n_6_2125), .A (n_6_1_224));
AOI222_X2 i_6_1_428 (.ZN (n_6_1_223), .A1 (n_6_1649), .A2 (drc_ipo_n26601), .B1 (n_6_1617)
    , .B2 (slo___n23215), .C1 (slo___n13169), .C2 (n_6_1_238));
INV_X2 i_6_1_427 (.ZN (n_6_2124), .A (n_6_1_223));
AOI222_X2 i_6_1_426 (.ZN (n_6_1_222), .A1 (n_6_1648), .A2 (drc_ipo_n26601), .B1 (n_6_1616)
    , .B2 (slo___n23215), .C1 (n_6_2155), .C2 (n_6_1_238));
INV_X2 i_6_1_425 (.ZN (n_6_2123), .A (n_6_1_222));
AOI222_X2 i_6_1_424 (.ZN (n_6_1_221), .A1 (n_6_1647), .A2 (drc_ipo_n26601), .B1 (n_6_1615)
    , .B2 (slo___n23215), .C1 (n_6_2154), .C2 (n_6_1_238));
INV_X2 i_6_1_423 (.ZN (n_6_2122), .A (n_6_1_221));
NAND2_X1 slo__sro_c21142 (.ZN (slo__sro_n18481), .A1 (CLOCK_sgo__n46934), .A2 (n_6_2736));
INV_X2 i_6_1_421 (.ZN (n_6_2121), .A (slo__sro_n18403));
AND2_X1 CLOCK_slo__sro_c54513 (.ZN (CLOCK_slo__sro_n49853), .A1 (n_6_90), .A2 (n_6_1_1079));
INV_X1 i_6_1_419 (.ZN (n_6_2120), .A (CLOCK_slo__sro_n52592));
AOI222_X2 i_6_1_418 (.ZN (n_6_1_218), .A1 (n_6_1644), .A2 (drc_ipo_n26601), .B1 (n_6_1612)
    , .B2 (slo___n23215), .C1 (n_6_2151), .C2 (n_6_1_238));
INV_X2 i_6_1_417 (.ZN (n_6_2119), .A (n_6_1_218));
AOI21_X1 CLOCK_slo__sro_c59417 (.ZN (CLOCK_slo__sro_n54100), .A (slo__sro_n4690), .B1 (n_6_1624), .B2 (slo___n23215));
AOI21_X4 CLOCK_sgo__sro_c51503 (.ZN (n_6_1_259), .A (CLOCK_sgo__sro_n47261), .B1 (n_6_1586), .B2 (slo___n23244));
AND2_X1 slo__sro_c17398 (.ZN (slo__sro_n15587), .A1 (n_6_2812), .A2 (n_6_1_973));
INV_X2 i_6_1_413 (.ZN (n_6_2117), .A (slo__sro_n15482));
AND2_X1 slo__sro_c6253 (.ZN (slo__sro_n5908), .A1 (n_6_2120), .A2 (n_6_1_203));
INV_X1 i_6_1_411 (.ZN (n_6_2116), .A (slo__sro_n5875));
NAND2_X1 slo__sro_c11661 (.ZN (slo__sro_n10771), .A1 (n_6_1817), .A2 (slo___n23226));
INV_X2 i_6_1_409 (.ZN (n_6_2115), .A (slo__sro_n10712));
INV_X1 CLOCK_slo__sro_c53347 (.ZN (CLOCK_slo__sro_n48815), .A (slo__sro_n20394));
INV_X2 i_6_1_407 (.ZN (n_6_2114), .A (n_6_1_213));
CLKBUF_X1 CLOCK_sgo__c52405 (.Z (CLOCK_sgo__n48008), .A (n_6_1_274));
INV_X2 i_6_1_405 (.ZN (n_6_2113), .A (n_6_1_212));
NAND2_X1 slo__sro_c22323 (.ZN (slo__sro_n19351), .A1 (n_6_2588), .A2 (n_6_1_728));
INV_X2 i_6_1_403 (.ZN (n_6_2112), .A (CLOCK_slo__sro_n51601));
AOI222_X1 i_6_1_402 (.ZN (n_6_1_210), .A1 (n_6_1636), .A2 (drc_ipo_n26601), .B1 (n_6_1604)
    , .B2 (slo___n23215), .C1 (n_6_2143), .C2 (n_6_1_238));
INV_X1 i_6_1_401 (.ZN (n_6_2111), .A (n_6_1_210));
AOI221_X2 slo__sro_c10133 (.ZN (slo__sro_n9429), .A (slo__sro_n9430), .B1 (n_6_988)
    , .B2 (slo___n23232), .C1 (n_6_1020), .C2 (slo___n23218));
INV_X4 i_6_1_399 (.ZN (n_6_2110), .A (slo__sro_n22024));
NAND2_X1 CLOCK_sgo__sro_c51750 (.ZN (CLOCK_sgo__sro_n47468), .A1 (CLOCK_sgo__sro_n47469), .A2 (CLOCK_sgo__sro_n47470));
INV_X2 i_6_1_397 (.ZN (n_6_2109), .A (n_6_1_208));
AOI222_X2 i_6_1_396 (.ZN (n_6_1_207), .A1 (n_6_1633), .A2 (drc_ipo_n26601), .B1 (n_6_1601)
    , .B2 (slo___n23215), .C1 (n_6_2140), .C2 (n_6_1_238));
INV_X2 i_6_1_395 (.ZN (n_6_2108), .A (n_6_1_207));
AOI222_X1 i_6_1_394 (.ZN (n_6_1_206), .A1 (n_6_1632), .A2 (drc_ipo_n26601), .B1 (n_6_1600)
    , .B2 (slo___n23215), .C1 (n_6_2139), .C2 (n_6_1_238));
INV_X1 i_6_1_393 (.ZN (n_6_2107), .A (n_6_1_206));
NOR2_X4 i_6_1_392 (.ZN (n_6_1_205), .A1 (n_6_1_1142), .A2 (Multiplicand[26]));
NOR2_X4 i_6_1_391 (.ZN (n_6_1_204), .A1 (Multiplicand[27]), .A2 (n_6_1_1141));
NOR2_X4 i_6_1_390 (.ZN (n_6_1_203), .A1 (slo___n23407), .A2 (slo___n23239));
AND2_X1 i_6_1_389 (.ZN (n_6_1_202), .A1 (n_6_2137), .A2 (n_6_1_203));
NAND2_X1 CLOCK_slo__sro_c56360 (.ZN (CLOCK_slo__sro_n51513), .A1 (n_6_2503), .A2 (n_6_1_623));
INV_X2 i_6_1_387 (.ZN (n_6_2106), .A (n_6_1_201));
AOI221_X2 i_6_1_386 (.ZN (n_6_1_200), .A (n_6_1_202), .B1 (n_6_1693), .B2 (n_6_1_204)
    , .C1 (n_6_1725), .C2 (slo___n23407));
INV_X2 i_6_1_385 (.ZN (n_6_2105), .A (n_6_1_200));
AOI21_X2 slo__sro_c6901 (.ZN (slo__sro_n6503), .A (slo__sro_n6504), .B1 (n_6_1273), .B2 (slo___n23274));
INV_X2 i_6_1_383 (.ZN (slo__n33292), .A (n_6_1_199));
AOI222_X2 slo__sro_c14593 (.ZN (slo__sro_n13262), .A1 (n_6_1845), .A2 (n_6_1_135)
    , .B1 (n_6_1813), .B2 (n_6_1_134), .C1 (slo__n17671), .C2 (n_6_1_133));
INV_X2 i_6_1_381 (.ZN (n_6_2103), .A (slo__sro_n13232));
NAND2_X1 slo__sro_c23313 (.ZN (slo__sro_n20262), .A1 (n_6_2496), .A2 (n_6_1_623));
INV_X2 i_6_1_379 (.ZN (n_6_2102), .A (CLOCK_slo__sro_n60309));
AND2_X1 slo__sro_c6871 (.ZN (slo__sro_n6480), .A1 (n_6_2161), .A2 (n_6_1_238));
INV_X2 i_6_1_377 (.ZN (n_6_2101), .A (n_6_1_196));
AOI222_X2 slo__sro_c37493 (.ZN (slo__sro_n33814), .A1 (n_6_1134), .A2 (slo___n23268)
    , .B1 (n_6_1102), .B2 (slo___n23277), .C1 (n_6_2401), .C2 (n_6_1_518));
INV_X2 i_6_1_375 (.ZN (n_6_2100), .A (slo__sro_n33595));
NAND2_X1 slo__sro_c33545 (.ZN (slo__sro_n30019), .A1 (n_6_816), .A2 (n_6_1_695));
INV_X1 i_6_1_373 (.ZN (slo___n18137), .A (slo__sro_n29857));
AOI222_X2 slo__sro_c15740 (.ZN (slo__sro_n14179), .A1 (n_6_1679), .A2 (n_6_1_204)
    , .B1 (n_6_1711), .B2 (slo___n23407), .C1 (n_6_2123), .C2 (n_6_1_203));
INV_X1 i_6_1_371 (.ZN (n_6_2098), .A (slo__sro_n14163));
AOI221_X2 slo__sro_c12820 (.ZN (slo__sro_n11754), .A (slo__sro_n11755), .B1 (n_6_1305)
    , .B2 (n_6_1_414), .C1 (n_6_1337), .C2 (slo___n43257));
INV_X2 i_6_1_369 (.ZN (spw__n69101), .A (slo__sro_n11728));
AOI222_X2 i_6_1_368 (.ZN (n_6_1_191), .A1 (n_6_1716), .A2 (slo___n23407), .B1 (n_6_1684)
    , .B2 (n_6_1_204), .C1 (n_6_2128), .C2 (n_6_1_203));
INV_X2 i_6_1_367 (.ZN (slo___n13213), .A (n_6_1_191));
INV_X1 slo__sro_c23686 (.ZN (slo__sro_n20615), .A (n_6_2847));
INV_X2 i_6_1_365 (.ZN (n_6_2095), .A (slo__sro_n20506));
NAND2_X1 slo__sro_c43067 (.ZN (slo__sro_n38916), .A1 (slo___n23359), .A2 (n_6_1232));
INV_X2 i_6_1_363 (.ZN (n_6_2094), .A (slo__sro_n14501));
AND2_X1 slo__sro_c11746 (.ZN (slo__sro_n10839), .A1 (n_6_2801), .A2 (n_6_1_973));
INV_X2 i_6_1_361 (.ZN (n_6_2093), .A (CLOCK_slo__sro_n60812));
NAND2_X1 slo__sro_c17276 (.ZN (slo__sro_n15472), .A1 (n_6_2109), .A2 (n_6_1_203));
INV_X1 i_6_1_359 (.ZN (n_6_2092), .A (n_6_1_187));
NAND2_X1 slo__sro_c15854 (.ZN (slo__sro_n14275), .A1 (CLOCK_sgo__n46945), .A2 (n_6_2876));
AND2_X2 slo__sro_c41457 (.ZN (slo__sro_n37539), .A1 (slo__sro_n37540), .A2 (slo__sro_n37541));
NAND2_X1 slo__sro_c14840 (.ZN (slo__sro_n13474), .A1 (slo__n32747), .A2 (n_6_1_378));
INV_X4 i_6_1_355 (.ZN (n_6_2090), .A (slo__sro_n13382));
NOR2_X1 slo__sro_c40161 (.ZN (slo__sro_n36417), .A1 (slo__sro_n36419), .A2 (slo__sro_n36418));
INV_X2 i_6_1_353 (.ZN (n_6_2089), .A (slo__sro_n36045));
NAND2_X1 slo__sro_c6312 (.ZN (slo__sro_n5965), .A1 (n_6_2614), .A2 (n_6_1_763));
INV_X2 i_6_1_351 (.ZN (n_6_2088), .A (slo__sro_n5907));
AND2_X1 slo__sro_c14939 (.ZN (slo__sro_n13545), .A1 (n_6_2746), .A2 (CLOCK_sgo__n46934));
INV_X2 i_6_1_349 (.ZN (n_6_2087), .A (n_6_1_182));
NAND2_X1 slo__sro_c16124 (.ZN (slo__sro_n14525), .A1 (slo__sro_n8872), .A2 (CLOCK_sgo__n46937));
INV_X2 i_6_1_347 (.ZN (n_6_2086), .A (slo__sro_n14441));
BUF_X32 drc_ipo_c29973 (.Z (drc_ipo_n26596), .A (slo__n3796));
INV_X1 i_6_1_345 (.ZN (n_6_2085), .A (n_6_1_180));
INV_X1 slo__sro_c34585 (.ZN (slo__sro_n30998), .A (slo__sro_n19776));
INV_X1 CLOCK_slo__sro_c56070 (.ZN (CLOCK_slo__sro_n51262), .A (slo__sro_n10370));
INV_X1 CLOCK_slo__sro_c59975 (.ZN (CLOCK_slo__sro_n54569), .A (slo__sro_n29226));
INV_X2 i_6_1_341 (.ZN (n_6_2083), .A (CLOCK_slo__sro_n54487));
AOI221_X2 CLOCK_slo__sro_c59891 (.ZN (CLOCK_slo__sro_n54487), .A (CLOCK_slo__sro_n54488)
    , .B1 (n_6_1671), .B2 (slo___n23239), .C1 (n_6_1703), .C2 (slo___n23407));
INV_X1 i_6_1_339 (.ZN (n_6_2082), .A (CLOCK_slo__sro_n54471));
NAND2_X1 slo__sro_c11660 (.ZN (slo__sro_n10772), .A1 (n_6_2071), .A2 (n_6_1_133));
INV_X1 i_6_1_337 (.ZN (n_6_2081), .A (slo__sro_n41478));
INV_X1 slo__sro_c10237 (.ZN (slo__sro_n9534), .A (slo__sro_n9535));
INV_X2 i_6_1_335 (.ZN (n_6_2080), .A (CLOCK_slo__sro_n48698));
INV_X1 slo__sro_c7051 (.ZN (slo__sro_n6652), .A (slo__sro_n6653));
INV_X2 i_6_1_333 (.ZN (n_6_2079), .A (CLOCK_slo__sro_n60762));
INV_X1 slo__sro_c33808 (.ZN (slo__sro_n30266), .A (slo__sro_n11035));
INV_X1 i_6_1_331 (.ZN (n_6_2078), .A (slo__sro_n30110));
NAND2_X1 slo__sro_c17292 (.ZN (slo__sro_n15485), .A1 (n_6_2149), .A2 (n_6_1_238));
INV_X2 i_6_1_329 (.ZN (n_6_2077), .A (n_6_1_172));
AOI222_X1 i_6_1_328 (.ZN (n_6_1_171), .A1 (n_6_1696), .A2 (slo___n23407), .B1 (n_6_1664)
    , .B2 (n_6_1_204), .C1 (n_6_2108), .C2 (n_6_1_203));
INV_X1 i_6_1_327 (.ZN (n_6_2076), .A (n_6_1_171));
NOR2_X2 i_6_1_326 (.ZN (n_6_1_170), .A1 (n_6_1_1143), .A2 (Multiplicand[27]));
NOR2_X4 i_6_1_325 (.ZN (n_6_1_169), .A1 (Multiplicand[28]), .A2 (n_6_1_1142));
NOR2_X4 i_6_1_324 (.ZN (n_6_1_168), .A1 (CLOCK_sgo__n48020), .A2 (slo___n23430));
AND2_X1 i_6_1_323 (.ZN (n_6_1_167), .A1 (n_6_2106), .A2 (n_6_1_168));
AOI222_X2 CLOCK_slo__sro_c58163 (.ZN (n_6_1_906), .A1 (n_6_320), .A2 (n_6_1_939), .B1 (n_6_352)
    , .B2 (n_6_1_940), .C1 (n_6_2759), .C2 (CLOCK_sgo__n46937));
INV_X4 i_6_1_321 (.ZN (n_6_2075), .A (n_6_1_166));
AOI221_X2 i_6_1_320 (.ZN (n_6_1_165), .A (n_6_1_167), .B1 (n_6_1757), .B2 (n_6_1_169)
    , .C1 (n_6_1789), .C2 (CLOCK_sgo__n48020));
INV_X1 i_6_1_319 (.ZN (n_6_2074), .A (n_6_1_165));
NAND2_X1 slo__sro_c14736 (.ZN (slo__sro_n13385), .A1 (n_6_2122), .A2 (n_6_1_203));
INV_X4 i_6_1_317 (.ZN (n_6_2073), .A (n_6_1_164));
AND2_X1 CLOCK_sgo__sro_c51900 (.ZN (CLOCK_sgo__sro_n47593), .A1 (n_6_2187), .A2 (n_6_1_273));
INV_X4 i_6_1_315 (.ZN (n_6_2072), .A (n_6_1_163));
AND2_X1 slo__sro_c35872 (.ZN (slo__sro_n32213), .A1 (n_6_1851), .A2 (n_6_1_135));
INV_X2 i_6_1_313 (.ZN (n_6_2071), .A (n_6_1_162));
AOI221_X1 slo__sro_c46789 (.ZN (slo__sro_n42331), .A (slo__sro_n42332), .B1 (n_6_742)
    , .B2 (n_6_1_730), .C1 (n_6_710), .C2 (n_6_1_729));
INV_X2 CLOCK_slo__c63328 (.ZN (CLOCK_slo__n57293), .A (slo__sro_n30110));
AOI21_X2 CLOCK_sgo__sro_c51479 (.ZN (n_6_1_155), .A (CLOCK_sgo__sro_n47244), .B1 (n_6_1747), .B2 (n_6_1_169));
INV_X2 i_6_1_309 (.ZN (n_6_2069), .A (n_6_1_160));
NAND2_X1 slo__sro_c14720 (.ZN (slo__sro_n13372), .A1 (n_6_1_168), .A2 (n_6_2105));
INV_X1 i_6_1_307 (.ZN (n_6_2068), .A (slo__sro_n13354));
AOI222_X2 i_6_1_306 (.ZN (n_6_1_158), .A1 (n_6_1782), .A2 (CLOCK_sgo__n48020), .B1 (n_6_1750)
    , .B2 (n_6_1_169), .C1 (n_6_2099), .C2 (n_6_1_168));
INV_X1 i_6_1_305 (.ZN (n_6_2067), .A (n_6_1_158));
AOI222_X1 CLOCK_slo__sro_c61778 (.ZN (n_6_1_994), .A1 (n_6_242), .A2 (n_6_1_1010)
    , .B1 (n_6_210), .B2 (n_6_1_1009), .C1 (n_6_2839), .C2 (CLOCK_sgo__n46950));
INV_X2 i_6_1_303 (.ZN (n_6_2066), .A (CLOCK_slo__sro_n51387));
NAND2_X1 slo__sro_c16536 (.ZN (slo__sro_n14856), .A1 (n_6_717), .A2 (n_6_1_729));
INV_X2 i_6_1_301 (.ZN (n_6_2065), .A (slo__sro_n27138));
INV_X1 i_6_1_299 (.ZN (n_6_2064), .A (n_6_1_155));
INV_X2 slo__c44046 (.ZN (slo__n39714), .A (slo__sro_n20506));
INV_X1 slo__c43729 (.ZN (slo__n39452), .A (slo__sro_n13461));
INV_X1 slo__c14627 (.ZN (slo__n13290), .A (n_6_1_69));
INV_X1 i_6_1_295 (.ZN (n_6_2062), .A (slo__sro_n13278));
INV_X1 slo__L1_c1_c39430 (.ZN (slo__n35732), .A (slo__n35733));
INV_X1 i_6_1_293 (.ZN (n_6_2061), .A (slo__sro_n14742));
AOI22_X4 slo__sro_c38440 (.ZN (slo__sro_n34792), .A1 (sgo__n1311), .A2 (sgo__n691)
    , .B1 (sgo__n1271), .B2 (sgo__n711));
INV_X1 i_6_1_291 (.ZN (n_6_2060), .A (slo__sro_n12647));
NAND2_X1 slo__sro_c17856 (.ZN (slo__sro_n15956), .A1 (n_6_1853), .A2 (n_6_1_135));
NAND2_X1 CLOCK_slo__sro_c53509 (.ZN (CLOCK_slo__sro_n48959), .A1 (n_6_1515), .A2 (slo___n23247));
NAND2_X4 CLOCK_slo__mro_c53132 (.ZN (slo__sro_n8603), .A1 (slo__sro_n8605), .A2 (slo__sro_n8604));
INV_X2 i_6_1_287 (.ZN (n_6_2058), .A (slo__sro_n15554));
AOI222_X2 i_6_1_286 (.ZN (n_6_1_148), .A1 (n_6_1772), .A2 (CLOCK_sgo__n48020), .B1 (n_6_1740)
    , .B2 (n_6_1_169), .C1 (n_6_2089), .C2 (n_6_1_168));
INV_X1 i_6_1_285 (.ZN (n_6_2057), .A (n_6_1_148));
NAND2_X4 slo__sro_c17500 (.ZN (slo__sro_n15669), .A1 (slo__sro_n15670), .A2 (slo__sro_n15671));
INV_X1 i_6_1_283 (.ZN (n_6_2056), .A (slo__sro_n15534));
AOI222_X2 i_6_1_282 (.ZN (n_6_1_146), .A1 (n_6_1770), .A2 (CLOCK_sgo__n48020), .B1 (n_6_1738)
    , .B2 (n_6_1_169), .C1 (n_6_2087), .C2 (n_6_1_168));
INV_X4 i_6_1_281 (.ZN (n_6_2055), .A (n_6_1_146));
AOI222_X2 i_6_1_280 (.ZN (n_6_1_145), .A1 (n_6_1769), .A2 (n_6_1_170), .B1 (n_6_1737)
    , .B2 (n_6_1_169), .C1 (n_6_2086), .C2 (n_6_1_168));
INV_X4 i_6_1_279 (.ZN (n_6_2054), .A (n_6_1_145));
NAND2_X1 slo__sro_c4888 (.ZN (slo__sro_n4674), .A1 (n_6_2861), .A2 (CLOCK_sgo__n46945));
INV_X1 i_6_1_277 (.ZN (n_6_2053), .A (slo__sro_n4615));
INV_X1 CLOCK_slo__sro_c67541 (.ZN (CLOCK_slo__sro_n60815), .A (slo__sro_n36567));
INV_X4 i_6_1_275 (.ZN (n_6_2052), .A (n_6_1_143));
NAND2_X1 CLOCK_slo__sro_c56310 (.ZN (CLOCK_slo__sro_n51473), .A1 (CLOCK_slo__sro_n51474), .A2 (CLOCK_slo__sro_n51475));
INV_X2 i_6_1_273 (.ZN (n_6_2051), .A (slo__sro_n39513));
AOI222_X2 i_6_1_272 (.ZN (n_6_1_141), .A1 (n_6_1765), .A2 (n_6_1_170), .B1 (n_6_1733)
    , .B2 (n_6_1_169), .C1 (n_6_2082), .C2 (n_6_1_168));
INV_X2 i_6_1_271 (.ZN (n_6_2050), .A (n_6_1_141));
NAND2_X1 slo__sro_c44165 (.ZN (slo__sro_n39795), .A1 (slo__sro_n39796), .A2 (slo__sro_n39797));
INV_X2 i_6_1_269 (.ZN (n_6_2049), .A (slo__sro_n39379));
AOI222_X2 i_6_1_268 (.ZN (n_6_1_139), .A1 (n_6_1763), .A2 (n_6_1_170), .B1 (n_6_1731)
    , .B2 (n_6_1_169), .C1 (n_6_2080), .C2 (n_6_1_168));
INV_X1 i_6_1_267 (.ZN (n_6_2048), .A (n_6_1_139));
AOI222_X2 i_6_1_266 (.ZN (n_6_1_138), .A1 (n_6_1762), .A2 (n_6_1_170), .B1 (n_6_1730)
    , .B2 (n_6_1_169), .C1 (n_6_2079), .C2 (n_6_1_168));
INV_X2 i_6_1_265 (.ZN (n_6_2047), .A (n_6_1_138));
AOI222_X2 i_6_1_264 (.ZN (n_6_1_137), .A1 (n_6_1761), .A2 (n_6_1_170), .B1 (n_6_1729)
    , .B2 (n_6_1_169), .C1 (n_6_2078), .C2 (n_6_1_168));
INV_X2 i_6_1_263 (.ZN (n_6_2046), .A (n_6_1_137));
AOI222_X1 i_6_1_262 (.ZN (n_6_1_136), .A1 (n_6_1760), .A2 (n_6_1_170), .B1 (n_6_1728)
    , .B2 (n_6_1_169), .C1 (n_6_2077), .C2 (n_6_1_168));
INV_X1 i_6_1_261 (.ZN (n_6_2045), .A (n_6_1_136));
NOR2_X4 i_6_1_260 (.ZN (n_6_1_135), .A1 (n_6_1_1144), .A2 (Multiplicand[28]));
NOR2_X4 i_6_1_259 (.ZN (n_6_1_134), .A1 (Multiplicand[29]), .A2 (n_6_1_1143));
NOR2_X4 i_6_1_258 (.ZN (n_6_1_133), .A1 (n_6_1_135), .A2 (n_6_1_134));
AND2_X1 i_6_1_257 (.ZN (n_6_1_132), .A1 (n_6_2075), .A2 (n_6_1_133));
AOI221_X2 i_6_1_256 (.ZN (n_6_1_131), .A (n_6_1_132), .B1 (n_6_1822), .B2 (spc__n66318)
    , .C1 (n_6_1854), .C2 (n_6_1_135));
INV_X2 i_6_1_255 (.ZN (n_6_2044), .A (n_6_1_131));
NAND2_X1 slo__sro_c18205 (.ZN (slo__sro_n16218), .A1 (n_6_2860), .A2 (CLOCK_sgo__n46945));
INV_X4 i_6_1_253 (.ZN (n_6_2043), .A (n_6_1_130));
AOI222_X2 i_6_1_252 (.ZN (n_6_1_129), .A1 (n_6_1852), .A2 (n_6_1_135), .B1 (n_6_1820)
    , .B2 (n_6_1_134), .C1 (n_6_2074), .C2 (n_6_1_133));
INV_X1 i_6_1_251 (.ZN (n_6_2042), .A (n_6_1_129));
INV_X1 slo__sro_c25890 (.ZN (slo__sro_n22624), .A (CLOCK_sgo__n46950));
INV_X1 i_6_1_249 (.ZN (n_6_2041), .A (slo__sro_n32212));
NAND2_X2 slo__sro_c31869 (.ZN (slo__sro_n28421), .A1 (n_6_968), .A2 (slo___n23232));
INV_X1 i_6_1_247 (.ZN (n_6_2040), .A (n_6_1_127));
INV_X2 i_6_1_245 (.ZN (n_6_2039), .A (slo__sro_n10769));
NAND2_X1 CLOCK_sgo__sro_c51346 (.ZN (CLOCK_sgo__sro_n47135), .A1 (n_6_1369), .A2 (n_6_1_379));
INV_X1 slo__c16346 (.ZN (slo__n14696), .A (slo__sro_n28523));
INV_X1 i_6_1_241 (.ZN (n_6_2037), .A (n_6_1_124));
NAND2_X1 slo__sro_c15724 (.ZN (slo__sro_n14166), .A1 (n_6_1_203), .A2 (n_6_2130));
INV_X1 i_6_1_239 (.ZN (n_6_2036), .A (n_6_1_123));
NAND2_X1 slo__sro_c14704 (.ZN (slo__sro_n13357), .A1 (n_6_2100), .A2 (n_6_1_168));
INV_X2 i_6_1_237 (.ZN (n_6_2035), .A (slo__sro_n13262));
AOI222_X2 i_6_1_236 (.ZN (n_6_1_121), .A1 (n_6_1844), .A2 (n_6_1_135), .B1 (n_6_1812)
    , .B2 (n_6_1_134), .C1 (n_6_2066), .C2 (n_6_1_133));
INV_X2 i_6_1_235 (.ZN (n_6_2034), .A (n_6_1_121));
AOI222_X2 i_6_1_234 (.ZN (n_6_1_120), .A1 (n_6_1843), .A2 (n_6_1_135), .B1 (n_6_1811)
    , .B2 (n_6_1_134), .C1 (n_6_2065), .C2 (n_6_1_133));
INV_X1 i_6_1_233 (.ZN (n_6_2033), .A (n_6_1_120));
AOI222_X2 CLOCK_slo__sro_c61291 (.ZN (CLOCK_slo__sro_n55687), .A1 (n_6_943), .A2 (n_6_1_625)
    , .B1 (n_6_911), .B2 (slo___n23367), .C1 (n_6_2495), .C2 (n_6_1_623));
INV_X1 i_6_1_231 (.ZN (n_6_2032), .A (CLOCK_slo__sro_n54789));
AOI222_X2 i_6_1_230 (.ZN (n_6_1_118), .A1 (n_6_1841), .A2 (n_6_1_135), .B1 (n_6_1809)
    , .B2 (n_6_1_134), .C1 (n_6_1_154), .C2 (n_6_1_133));
INV_X2 i_6_1_229 (.ZN (n_6_2031), .A (n_6_1_118));
AOI222_X2 i_6_1_228 (.ZN (n_6_1_117), .A1 (n_6_1840), .A2 (n_6_1_135), .B1 (n_6_1808)
    , .B2 (slo___n43254), .C1 (n_6_2062), .C2 (n_6_1_133));
INV_X1 i_6_1_227 (.ZN (slo___n15411), .A (n_6_1_117));
AOI222_X2 slo__sro_c17363 (.ZN (slo__sro_n15554), .A1 (n_6_1741), .A2 (n_6_1_169)
    , .B1 (n_6_1773), .B2 (CLOCK_sgo__n48020), .C1 (n_6_2090), .C2 (n_6_1_168));
BUF_X1 slo__L3_c3_c30024 (.Z (slo__n26654), .A (n_6_8));
AOI222_X2 i_6_1_224 (.ZN (n_6_1_115), .A1 (n_6_1838), .A2 (n_6_1_135), .B1 (n_6_1806)
    , .B2 (n_6_1_134), .C1 (n_6_2060), .C2 (n_6_1_133));
NAND2_X1 CLOCK_sgo__sro_c51749 (.ZN (CLOCK_sgo__sro_n47469), .A1 (n_6_1755), .A2 (n_6_1_169));
AOI222_X2 slo__sro_c7239 (.ZN (slo__sro_n6817), .A1 (n_6_1186), .A2 (slo___n23466)
    , .B1 (n_6_1154), .B2 (slo___n23364), .C1 (slo___n17582), .C2 (n_6_1_483));
INV_X1 i_6_1_221 (.ZN (n_6_2027), .A (slo__sro_n6737));
AOI221_X2 slo__sro_c6872 (.ZN (slo__sro_n6479), .A (slo__sro_n6480), .B1 (n_6_1622)
    , .B2 (slo___n23215), .C1 (n_6_1654), .C2 (drc_ipo_n26601));
INV_X2 i_6_1_219 (.ZN (n_6_2026), .A (slo__sro_n6366));
INV_X1 CLOCK_slo__sro_c53581 (.ZN (CLOCK_slo__sro_n49025), .A (slo__sro_n40292));
INV_X2 i_6_1_217 (.ZN (n_6_2025), .A (n_6_1_112));
NOR2_X1 slo__sro_c11192 (.ZN (slo__sro_n10378), .A1 (slo__sro_n10380), .A2 (slo__sro_n10379));
INV_X2 i_6_1_215 (.ZN (n_6_2024), .A (slo__sro_n10311));
AND2_X1 slo__sro_c11594 (.ZN (slo__sro_n10713), .A1 (n_6_2147), .A2 (n_6_1_238));
INV_X2 i_6_1_213 (.ZN (n_6_2023), .A (CLOCK_slo__sro_n60603));
AOI221_X2 CLOCK_sgo__sro_c51901 (.ZN (spt__n66402), .A (CLOCK_sgo__sro_n47593), .B1 (n_6_1553)
    , .B2 (n_6_1_274), .C1 (n_6_1585), .C2 (slo___n23244));
INV_X1 i_6_1_211 (.ZN (n_6_2022), .A (n_6_1_109));
AOI222_X2 CLOCK_slo__sro_c59754 (.ZN (n_6_1_1053), .A1 (n_6_103), .A2 (n_6_1_1080)
    , .B1 (n_6_71), .B2 (n_6_1_1079), .C1 (slo__n12005), .C2 (slo__n13799));
INV_X1 i_6_1_209 (.ZN (n_6_2021), .A (CLOCK_slo__sro_n54312));
AOI222_X2 i_6_1_208 (.ZN (spw__n67541), .A1 (n_6_1830), .A2 (n_6_1_135), .B1 (n_6_1798)
    , .B2 (n_6_1_134), .C1 (n_6_2052), .C2 (n_6_1_133));
AOI221_X2 slo__sro_c32553 (.ZN (slo__sro_n29067), .A (slo__sro_n29068), .B1 (n_6_1796)
    , .B2 (n_6_1_134), .C1 (n_6_1828), .C2 (slo___n23404));
NAND2_X1 CLOCK_slo__sro_c68792 (.ZN (CLOCK_slo__sro_n61963), .A1 (n_6_2372), .A2 (n_6_1_483));
INV_X2 i_6_1_205 (.ZN (n_6_2019), .A (CLOCK_slo__sro_n61783));
NOR2_X1 slo__sro_c32724 (.ZN (slo__sro_n29226), .A1 (slo__sro_n29228), .A2 (slo__sro_n29227));
INV_X2 i_6_1_203 (.ZN (n_6_2018), .A (slo__sro_n29067));
INV_X1 slo__sro_c32552 (.ZN (slo__sro_n29068), .A (slo__sro_n29069));
INV_X2 i_6_1_201 (.ZN (n_6_2017), .A (slo__sro_n29017));
INV_X1 CLOCK_slo__sro_c60516 (.ZN (CLOCK_slo__sro_n55023), .A (slo__sro_n6283));
INV_X2 i_6_1_199 (.ZN (n_6_2016), .A (n_6_1_103));
AOI222_X2 i_6_1_198 (.ZN (n_6_1_102), .A1 (n_6_1825), .A2 (slo___n23404), .B1 (n_6_1793)
    , .B2 (n_6_1_134), .C1 (n_6_2047), .C2 (n_6_1_133));
INV_X2 i_6_1_197 (.ZN (n_6_2015), .A (n_6_1_102));
AOI222_X1 i_6_1_196 (.ZN (n_6_1_101), .A1 (n_6_1824), .A2 (slo___n23404), .B1 (n_6_1792)
    , .B2 (n_6_1_134), .C1 (n_6_2046), .C2 (n_6_1_133));
INV_X1 i_6_1_195 (.ZN (n_6_2014), .A (n_6_1_101));
NOR2_X1 i_6_1_194 (.ZN (CLOCK_slo__n60586), .A1 (n_6_1_1145), .A2 (Multiplicand[29]));
NOR2_X2 i_6_1_193 (.ZN (n_6_1_99), .A1 (Multiplicand[30]), .A2 (n_6_1_1144));
NOR2_X4 i_6_1_192 (.ZN (n_6_1_98), .A1 (n_6_1_100), .A2 (CLOCK_sgo__n48011));
AND2_X1 i_6_1_191 (.ZN (n_6_1_97), .A1 (n_6_2044), .A2 (n_6_1_98));
AOI221_X2 i_6_1_190 (.ZN (n_6_1_96), .A (n_6_1_97), .B1 (n_6_1886), .B2 (n_6_1_99)
    , .C1 (n_6_1918), .C2 (slo___n43247));
INV_X1 i_6_1_189 (.ZN (n_6_2013), .A (n_6_1_96));
AOI221_X2 i_6_1_188 (.ZN (n_6_1_95), .A (n_6_1_97), .B1 (n_6_1885), .B2 (n_6_1_99)
    , .C1 (n_6_1917), .C2 (n_6_1_100));
INV_X4 i_6_1_187 (.ZN (n_6_2012), .A (n_6_1_95));
AOI222_X2 i_6_1_186 (.ZN (n_6_1_94), .A1 (n_6_1916), .A2 (slo___n23235), .B1 (n_6_1884)
    , .B2 (slo___n23221), .C1 (n_6_2043), .C2 (n_6_1_98));
INV_X2 i_6_1_185 (.ZN (n_6_2011), .A (n_6_1_94));
NAND2_X1 CLOCK_slo__sro_c65159 (.ZN (CLOCK_slo__sro_n58710), .A1 (n_6_1626), .A2 (slo___n23215));
INV_X2 i_6_1_183 (.ZN (n_6_2010), .A (n_6_1_93));
NAND2_X1 slo__sro_c30754 (.ZN (slo__sro_n27361), .A1 (n_6_793), .A2 (n_6_1_694));
INV_X4 i_6_1_181 (.ZN (n_6_2009), .A (slo__sro_n34317));
AND2_X1 slo__sro_c10132 (.ZN (slo__sro_n9430), .A1 (n_6_2477), .A2 (n_6_1_588));
NAND2_X1 slo__sro_c30903 (.ZN (slo__sro_n27501), .A1 (n_6_1_995), .A2 (n_6_1_973));
NAND2_X1 CLOCK_slo__sro_c68794 (.ZN (CLOCK_slo__sro_n61961), .A1 (CLOCK_slo__sro_n61962), .A2 (CLOCK_slo__sro_n61963));
INV_X2 i_6_1_177 (.ZN (n_6_2007), .A (n_6_1_90));
CLKBUF_X1 slo__L3_c3_c43528 (.Z (n_6_1_154), .A (slo__n39284));
INV_X2 i_6_1_175 (.ZN (n_6_2006), .A (slo__sro_n39249));
INV_X2 i_6_1_173 (.ZN (slo__n40097), .A (n_6_1_88));
AOI222_X2 i_6_1_172 (.ZN (n_6_1_87), .A1 (n_6_1909), .A2 (n_6_1_100), .B1 (n_6_1877)
    , .B2 (CLOCK_sgo__n48011), .C1 (n_6_2036), .C2 (n_6_1_98));
INV_X2 i_6_1_171 (.ZN (n_6_2004), .A (n_6_1_87));
AOI222_X1 i_6_1_170 (.ZN (n_6_1_86), .A1 (n_6_1908), .A2 (n_6_1_100), .B1 (n_6_1876)
    , .B2 (CLOCK_sgo__n48011), .C1 (n_6_2035), .C2 (n_6_1_98));
INV_X2 i_6_1_169 (.ZN (n_6_2003), .A (n_6_1_86));
AOI222_X1 i_6_1_168 (.ZN (n_6_1_85), .A1 (n_6_1907), .A2 (n_6_1_100), .B1 (n_6_1875)
    , .B2 (CLOCK_sgo__n48011), .C1 (n_6_2034), .C2 (n_6_1_98));
INV_X2 i_6_1_167 (.ZN (n_6_2002), .A (n_6_1_85));
AOI222_X1 i_6_1_166 (.ZN (n_6_1_84), .A1 (n_6_1906), .A2 (n_6_1_100), .B1 (n_6_1874)
    , .B2 (CLOCK_sgo__n48011), .C1 (n_6_2033), .C2 (n_6_1_98));
INV_X1 i_6_1_165 (.ZN (n_6_2001), .A (n_6_1_84));
AOI222_X1 i_6_1_164 (.ZN (n_6_1_83), .A1 (n_6_1905), .A2 (n_6_1_100), .B1 (n_6_1873)
    , .B2 (CLOCK_sgo__n48011), .C1 (n_6_2032), .C2 (n_6_1_98));
INV_X1 i_6_1_163 (.ZN (n_6_2000), .A (n_6_1_83));
AOI222_X1 i_6_1_162 (.ZN (n_6_1_82), .A1 (n_6_1904), .A2 (n_6_1_100), .B1 (n_6_1872)
    , .B2 (CLOCK_sgo__n48011), .C1 (n_6_2031), .C2 (n_6_1_98));
INV_X1 i_6_1_161 (.ZN (n_6_1999), .A (n_6_1_82));
AOI222_X1 i_6_1_160 (.ZN (n_6_1_81), .A1 (n_6_1903), .A2 (n_6_1_100), .B1 (n_6_1871)
    , .B2 (CLOCK_sgo__n48011), .C1 (slo___n15411), .C2 (n_6_1_98));
INV_X1 i_6_1_159 (.ZN (n_6_1998), .A (n_6_1_81));
NAND2_X1 CLOCK_slo__sro_c56762 (.ZN (CLOCK_slo__sro_n51853), .A1 (n_6_1572), .A2 (slo___n23244));
INV_X1 i_6_1_157 (.ZN (n_6_1997), .A (CLOCK_slo__sro_n51773));
AOI222_X1 i_6_1_156 (.ZN (n_6_1_79), .A1 (n_6_1901), .A2 (n_6_1_100), .B1 (n_6_1869)
    , .B2 (CLOCK_sgo__n48011), .C1 (CLOCK_opt_ipo_n45742), .C2 (n_6_1_98));
INV_X1 i_6_1_155 (.ZN (n_6_1996), .A (n_6_1_79));
AOI222_X1 i_6_1_154 (.ZN (n_6_1_78), .A1 (n_6_1900), .A2 (n_6_1_100), .B1 (n_6_1868)
    , .B2 (CLOCK_sgo__n48011), .C1 (opt_ipo_n24196), .C2 (n_6_1_98));
INV_X1 i_6_1_153 (.ZN (n_6_1995), .A (n_6_1_78));
AOI222_X2 i_6_1_152 (.ZN (n_6_1_77), .A1 (n_6_1899), .A2 (n_6_1_100), .B1 (n_6_1867)
    , .B2 (CLOCK_sgo__n48011), .C1 (n_6_2026), .C2 (n_6_1_98));
INV_X1 i_6_1_151 (.ZN (n_6_1994), .A (n_6_1_77));
INV_X2 CLOCK_slo__c63265 (.ZN (CLOCK_slo__n57242), .A (slo__sro_n32212));
INV_X2 i_6_1_149 (.ZN (spw__n68268), .A (CLOCK_slo__sro_n57132));
AOI221_X2 CLOCK_slo__sro_c72495 (.ZN (n_6_1_1040), .A (n_6_1_1042), .B1 (n_6_157)
    , .B2 (n_6_1_1044), .C1 (n_6_189), .C2 (n_6_1_1045));
INV_X1 i_6_1_147 (.ZN (n_6_1992), .A (slo__sro_n39363));
AOI222_X2 slo__sro_c11344 (.ZN (n_6_1_68), .A1 (n_6_1858), .A2 (n_6_1_99), .B1 (n_6_1890)
    , .B2 (n_6_1_100), .C1 (n_6_2017), .C2 (n_6_1_98));
AOI222_X2 slo__sro_c43644 (.ZN (slo__sro_n39379), .A1 (n_6_1732), .A2 (n_6_1_169)
    , .B1 (n_6_1764), .B2 (n_6_1_170), .C1 (n_6_2081), .C2 (n_6_1_168));
INV_X1 i_6_1_143 (.ZN (n_6_1990), .A (n_6_1_73));
NAND2_X1 slo__sro_c12636 (.ZN (slo__sro_n11596), .A1 (n_6_1308), .A2 (n_6_1_414));
INV_X1 i_6_1_141 (.ZN (n_6_1989), .A (slo__sro_n11496));
AOI222_X2 slo__sro_c6784 (.ZN (n_6_1_196), .A1 (n_6_1721), .A2 (slo___n23407), .B1 (n_6_1689)
    , .B2 (n_6_1_204), .C1 (n_6_2133), .C2 (n_6_1_203));
INV_X2 i_6_1_139 (.ZN (n_6_1988), .A (CLOCK_slo__sro_n64581));
AOI222_X2 i_6_1_138 (.ZN (n_6_1_70), .A1 (n_6_1892), .A2 (n_6_1_100), .B1 (n_6_1860)
    , .B2 (n_6_1_99), .C1 (n_6_2019), .C2 (n_6_1_98));
INV_X1 i_6_1_137 (.ZN (n_6_1987), .A (n_6_1_70));
AOI222_X2 i_6_1_136 (.ZN (n_6_1_69), .A1 (n_6_1891), .A2 (n_6_1_100), .B1 (n_6_1859)
    , .B2 (n_6_1_99), .C1 (n_6_2018), .C2 (n_6_1_98));
INV_X1 i_6_1_135 (.ZN (n_6_1986), .A (n_6_1_69));
NAND2_X1 slo__sro_c40638 (.ZN (slo__sro_n36836), .A1 (n_6_1116), .A2 (slo___n23277));
INV_X2 i_6_1_133 (.ZN (n_6_1985), .A (n_6_1_68));
AOI222_X2 i_6_1_132 (.ZN (n_6_1_67), .A1 (n_6_1889), .A2 (n_6_1_100), .B1 (n_6_1857)
    , .B2 (n_6_1_99), .C1 (n_6_2016), .C2 (n_6_1_98));
INV_X2 i_6_1_131 (.ZN (n_6_1984), .A (n_6_1_67));
AOI222_X1 i_6_1_130 (.ZN (n_6_1_66), .A1 (n_6_1888), .A2 (n_6_1_100), .B1 (n_6_1856)
    , .B2 (n_6_1_99), .C1 (n_6_2015), .C2 (n_6_1_98));
INV_X1 i_6_1_129 (.ZN (n_6_1983), .A (n_6_1_66));
AND2_X4 i_6_1_128 (.ZN (n_6_1_65), .A1 (Multiplicand[31]), .A2 (n_6_1_1145));
NOR2_X4 i_6_1_127 (.ZN (n_6_1_64), .A1 (Multiplicand[31]), .A2 (n_6_1_1145));
NOR2_X4 i_6_1_126 (.ZN (n_6_1_63), .A1 (n_6_1_65), .A2 (n_6_1_64));
AND2_X1 i_6_1_125 (.ZN (n_6_1_62), .A1 (n_6_2013), .A2 (n_6_1_63));
AOI21_X4 slo__sro_c2007 (.ZN (slo__sro_n2106), .A (slo__sro_n2107), .B1 (n_6_38), .B2 (n_6_1_1114));
NAND2_X1 CLOCK_slo__sro_c68772 (.ZN (CLOCK_slo__sro_n61943), .A1 (CLOCK_slo__sro_n61944), .A2 (CLOCK_slo__sro_n61945));
INV_X1 slo__mro_c36953 (.ZN (slo__mro_n33302), .A (hfn_ipo_n35));
NAND2_X2 slo__sro_c37268 (.ZN (slo__sro_n33597), .A1 (n_6_1688), .A2 (n_6_1_204));
NAND2_X2 slo__sro_c37269 (.ZN (slo__sro_n33596), .A1 (slo__sro_n33597), .A2 (slo__sro_n33598));
AOI222_X2 i_6_1_118 (.ZN (n_6_1_58), .A1 (n_6_1979), .A2 (n_6_1_65), .B1 (n_6_1947)
    , .B2 (n_6_1_64), .C1 (slo__n13053), .C2 (n_6_1_63));
NAND2_X1 CLOCK_slo__sro_c56674 (.ZN (CLOCK_slo__sro_n51775), .A1 (n_6_1902), .A2 (n_6_1_100));
INV_X8 CLOCK_slo__c55144 (.ZN (CLOCK_slo__n50421), .A (CLOCK_slo__n50420));
AOI222_X1 slo__sro_c14326 (.ZN (slo__sro_n13037), .A1 (n_6_1978), .A2 (n_6_1_65), .B1 (n_6_1946)
    , .B2 (n_6_1_64), .C1 (n_6_2010), .C2 (n_6_1_63));
INV_X1 i_6_1_113 (.ZN (n_57), .A (slo__sro_n13019));
AOI222_X2 i_6_1_112 (.ZN (n_6_1_55), .A1 (n_6_1976), .A2 (n_6_1_65), .B1 (n_6_1944)
    , .B2 (n_6_1_64), .C1 (slo__n27410), .C2 (n_6_1_63));
INV_X1 i_6_1_111 (.ZN (n_56), .A (n_6_1_55));
AOI222_X1 i_6_1_110 (.ZN (n_6_1_54), .A1 (n_6_1975), .A2 (n_6_1_65), .B1 (n_6_1943)
    , .B2 (n_6_1_64), .C1 (n_6_2007), .C2 (n_6_1_63));
INV_X1 i_6_1_109 (.ZN (n_55), .A (n_6_1_54));
OR2_X4 CLOCK_slo__c62386 (.ZN (slo__sro_n8872), .A1 (slo__sro_n8873), .A2 (CLOCK_slo__sro_n56306));
INV_X1 i_6_1_107 (.ZN (n_54), .A (n_6_1_53));
AOI222_X1 i_6_1_106 (.ZN (CLOCK_slo__n54298), .A1 (n_6_1973), .A2 (n_6_1_65), .B1 (n_6_1941)
    , .B2 (n_6_1_64), .C1 (slo__n40097), .C2 (n_6_1_63));
INV_X2 CLOCK_slo__c60093 (.ZN (CLOCK_slo__n54661), .A (n_6_1_436));
AOI222_X1 i_6_1_104 (.ZN (n_6_1_51), .A1 (n_6_1972), .A2 (n_6_1_65), .B1 (n_6_1940)
    , .B2 (n_6_1_64), .C1 (n_6_2004), .C2 (n_6_1_63));
INV_X1 i_6_1_103 (.ZN (n_52), .A (n_6_1_51));
AOI222_X1 i_6_1_102 (.ZN (n_6_1_50), .A1 (n_6_1971), .A2 (n_6_1_65), .B1 (n_6_1939)
    , .B2 (n_6_1_64), .C1 (n_6_2003), .C2 (n_6_1_63));
INV_X1 i_6_1_101 (.ZN (n_51), .A (n_6_1_50));
AOI222_X1 i_6_1_100 (.ZN (n_6_1_49), .A1 (n_6_1970), .A2 (n_6_1_65), .B1 (n_6_1938)
    , .B2 (n_6_1_64), .C1 (n_6_2002), .C2 (n_6_1_63));
INV_X1 i_6_1_99 (.ZN (n_50), .A (n_6_1_49));
AOI222_X1 i_6_1_98 (.ZN (n_6_1_48), .A1 (n_6_1969), .A2 (n_6_1_65), .B1 (n_6_1937)
    , .B2 (n_6_1_64), .C1 (n_6_2001), .C2 (n_6_1_63));
INV_X1 i_6_1_97 (.ZN (n_49), .A (n_6_1_48));
AOI222_X1 i_6_1_96 (.ZN (spt__n66349), .A1 (n_6_1968), .A2 (n_6_1_65), .B1 (n_6_1936)
    , .B2 (n_6_1_64), .C1 (n_6_2000), .C2 (n_6_1_63));
INV_X1 i_6_1_95 (.ZN (n_48), .A (n_6_1_47));
AOI222_X1 i_6_1_94 (.ZN (n_6_1_46), .A1 (n_6_1967), .A2 (n_6_1_65), .B1 (n_6_1935)
    , .B2 (n_6_1_64), .C1 (n_6_1999), .C2 (n_6_1_63));
INV_X1 i_6_1_93 (.ZN (n_47), .A (n_6_1_46));
AOI222_X1 i_6_1_92 (.ZN (n_6_1_45), .A1 (n_6_1966), .A2 (n_6_1_65), .B1 (n_6_1934)
    , .B2 (n_6_1_64), .C1 (n_6_1998), .C2 (n_6_1_63));
INV_X1 i_6_1_91 (.ZN (n_46), .A (n_6_1_45));
AOI222_X1 i_6_1_90 (.ZN (n_6_1_44), .A1 (n_6_1965), .A2 (n_6_1_65), .B1 (n_6_1933)
    , .B2 (n_6_1_64), .C1 (n_6_1997), .C2 (n_6_1_63));
INV_X1 i_6_1_89 (.ZN (n_45), .A (n_6_1_44));
AOI222_X1 i_6_1_88 (.ZN (n_6_1_43), .A1 (n_6_1964), .A2 (n_6_1_65), .B1 (n_6_1932)
    , .B2 (n_6_1_64), .C1 (n_6_1996), .C2 (n_6_1_63));
INV_X1 i_6_1_87 (.ZN (n_44), .A (n_6_1_43));
AOI222_X1 i_6_1_86 (.ZN (n_6_1_42), .A1 (n_6_1963), .A2 (n_6_1_65), .B1 (n_6_1931)
    , .B2 (n_6_1_64), .C1 (n_6_1995), .C2 (n_6_1_63));
INV_X1 i_6_1_85 (.ZN (n_43), .A (n_6_1_42));
AOI222_X1 i_6_1_84 (.ZN (n_6_1_41), .A1 (n_6_1962), .A2 (n_6_1_65), .B1 (n_6_1930)
    , .B2 (n_6_1_64), .C1 (n_6_1994), .C2 (n_6_1_63));
INV_X1 i_6_1_83 (.ZN (n_42), .A (n_6_1_41));
AOI222_X1 i_6_1_82 (.ZN (n_6_1_40), .A1 (n_6_1961), .A2 (n_6_1_65), .B1 (n_6_1929)
    , .B2 (n_6_1_64), .C1 (n_6_1993), .C2 (n_6_1_63));
INV_X1 i_6_1_81 (.ZN (n_41), .A (n_6_1_40));
AOI222_X1 i_6_1_80 (.ZN (n_6_1_39), .A1 (n_6_1960), .A2 (n_6_1_65), .B1 (n_6_1928)
    , .B2 (n_6_1_64), .C1 (n_6_1992), .C2 (n_6_1_63));
INV_X1 i_6_1_79 (.ZN (n_40), .A (n_6_1_39));
AOI222_X1 i_6_1_78 (.ZN (n_6_1_38), .A1 (n_6_1959), .A2 (n_6_1_65), .B1 (n_6_1927)
    , .B2 (n_6_1_64), .C1 (n_6_1_74), .C2 (n_6_1_63));
INV_X1 i_6_1_77 (.ZN (n_39), .A (n_6_1_38));
AOI222_X1 i_6_1_76 (.ZN (n_6_1_37), .A1 (n_6_1958), .A2 (n_6_1_65), .B1 (n_6_1926)
    , .B2 (n_6_1_64), .C1 (n_6_1990), .C2 (n_6_1_63));
INV_X1 i_6_1_75 (.ZN (n_38), .A (n_6_1_37));
AOI222_X1 i_6_1_74 (.ZN (n_6_1_36), .A1 (n_6_1957), .A2 (n_6_1_65), .B1 (n_6_1925)
    , .B2 (n_6_1_64), .C1 (n_6_1989), .C2 (n_6_1_63));
INV_X1 i_6_1_73 (.ZN (n_37), .A (n_6_1_36));
AOI222_X1 i_6_1_72 (.ZN (n_6_1_35), .A1 (n_6_1956), .A2 (n_6_1_65), .B1 (n_6_1924)
    , .B2 (n_6_1_64), .C1 (n_6_1988), .C2 (n_6_1_63));
INV_X1 i_6_1_71 (.ZN (n_36), .A (n_6_1_35));
AOI222_X1 i_6_1_70 (.ZN (n_6_1_34), .A1 (n_6_1955), .A2 (n_6_1_65), .B1 (n_6_1923)
    , .B2 (n_6_1_64), .C1 (n_6_1987), .C2 (n_6_1_63));
INV_X1 i_6_1_69 (.ZN (n_35), .A (n_6_1_34));
AOI222_X1 i_6_1_68 (.ZN (n_6_1_33), .A1 (n_6_1954), .A2 (n_6_1_65), .B1 (n_6_1922)
    , .B2 (n_6_1_64), .C1 (n_6_1986), .C2 (n_6_1_63));
INV_X1 i_6_1_67 (.ZN (n_34), .A (n_6_1_33));
AOI222_X1 i_6_1_66 (.ZN (n_6_1_32), .A1 (n_6_1953), .A2 (n_6_1_65), .B1 (n_6_1921)
    , .B2 (n_6_1_64), .C1 (n_6_1985), .C2 (n_6_1_63));
INV_X1 i_6_1_65 (.ZN (n_33), .A (n_6_1_32));
AOI222_X1 i_6_1_64 (.ZN (n_6_1_31), .A1 (n_6_1952), .A2 (n_6_1_65), .B1 (n_6_1920)
    , .B2 (n_6_1_64), .C1 (n_6_1984), .C2 (n_6_1_63));
INV_X1 i_6_1_63 (.ZN (n_32), .A (n_6_1_31));
AOI222_X1 i_6_1_62 (.ZN (n_6_1_30), .A1 (n_6_1951), .A2 (n_6_1_65), .B1 (n_6_1919)
    , .B2 (n_6_1_64), .C1 (n_6_1983), .C2 (n_6_1_63));
INV_X1 i_6_1_61 (.ZN (n_31), .A (n_6_1_30));
AOI222_X2 i_6_1_60 (.ZN (n_6_1_29), .A1 (n_6_1887), .A2 (n_6_1_100), .B1 (n_6_1855)
    , .B2 (n_6_1_99), .C1 (n_6_2014), .C2 (n_6_1_98));
INV_X1 i_6_1_59 (.ZN (n_30), .A (n_6_1_29));
AOI222_X1 i_6_1_58 (.ZN (n_6_1_28), .A1 (n_6_1823), .A2 (slo___n23404), .B1 (n_6_1791)
    , .B2 (n_6_1_134), .C1 (n_6_2045), .C2 (n_6_1_133));
INV_X1 i_6_1_57 (.ZN (n_29), .A (n_6_1_28));
AOI222_X1 i_6_1_56 (.ZN (n_6_1_27), .A1 (n_6_1759), .A2 (CLOCK_sgo__n48020), .B1 (n_6_1727)
    , .B2 (n_6_1_169), .C1 (n_6_2076), .C2 (n_6_1_168));
INV_X1 i_6_1_55 (.ZN (n_28), .A (n_6_1_27));
AOI222_X1 i_6_1_54 (.ZN (n_6_1_26), .A1 (n_6_1695), .A2 (slo___n23407), .B1 (n_6_1663)
    , .B2 (n_6_1_204), .C1 (n_6_2107), .C2 (n_6_1_203));
INV_X1 i_6_1_53 (.ZN (n_27), .A (n_6_1_26));
AOI222_X1 i_6_1_52 (.ZN (n_6_1_25), .A1 (n_6_1631), .A2 (drc_ipo_n26601), .B1 (n_6_1599)
    , .B2 (slo___n23215), .C1 (n_6_2138), .C2 (n_6_1_238));
INV_X1 i_6_1_51 (.ZN (n_26), .A (n_6_1_25));
AOI222_X1 i_6_1_50 (.ZN (n_6_1_24), .A1 (n_6_1567), .A2 (slo___n23244), .B1 (n_6_1535)
    , .B2 (n_6_1_274), .C1 (n_6_2169), .C2 (n_6_1_273));
INV_X1 i_6_1_49 (.ZN (n_25), .A (n_6_1_24));
AOI222_X1 i_6_1_48 (.ZN (n_6_1_23), .A1 (n_6_1503), .A2 (slo___n23247), .B1 (n_6_1471)
    , .B2 (n_6_1_309), .C1 (n_6_2200), .C2 (n_6_1_308));
INV_X1 i_6_1_47 (.ZN (n_24), .A (n_6_1_23));
AOI222_X1 i_6_1_46 (.ZN (n_6_1_22), .A1 (n_6_1439), .A2 (n_6_1_345), .B1 (n_6_1407)
    , .B2 (slo___n23229), .C1 (n_6_2231), .C2 (n_6_1_343));
INV_X1 i_6_1_45 (.ZN (n_23), .A (n_6_1_22));
AOI222_X1 i_6_1_44 (.ZN (n_6_1_21), .A1 (n_6_1375), .A2 (n_6_1_380), .B1 (n_6_1343)
    , .B2 (n_6_1_379), .C1 (n_6_2262), .C2 (n_6_1_378));
INV_X1 i_6_1_43 (.ZN (n_22), .A (n_6_1_21));
AOI222_X1 i_6_1_42 (.ZN (n_6_1_20), .A1 (n_6_1279), .A2 (n_6_1_414), .B1 (n_6_1311)
    , .B2 (slo___n43257), .C1 (n_6_2293), .C2 (n_6_1_413));
INV_X1 i_6_1_41 (.ZN (n_21), .A (n_6_1_20));
AOI222_X1 i_6_1_40 (.ZN (n_6_1_19), .A1 (n_6_1215), .A2 (slo___n23359), .B1 (n_6_1247)
    , .B2 (slo___n23274), .C1 (n_6_2324), .C2 (n_6_1_448));
INV_X1 i_6_1_39 (.ZN (n_20), .A (n_6_1_19));
AOI222_X1 i_6_1_38 (.ZN (n_6_1_18), .A1 (n_6_1151), .A2 (slo___n23364), .B1 (n_6_1183)
    , .B2 (slo___n23466), .C1 (n_6_2355), .C2 (n_6_1_483));
INV_X1 i_6_1_37 (.ZN (n_19), .A (n_6_1_18));
AOI222_X1 i_6_1_36 (.ZN (n_6_1_17), .A1 (n_6_1087), .A2 (slo___n23277), .B1 (n_6_1119)
    , .B2 (slo___n23268), .C1 (n_6_2386), .C2 (n_6_1_518));
INV_X1 i_6_1_35 (.ZN (n_18), .A (n_6_1_17));
AOI222_X1 i_6_1_34 (.ZN (n_6_1_16), .A1 (n_6_1023), .A2 (slo___n23353), .B1 (n_6_1055)
    , .B2 (slo___n23457), .C1 (n_6_2417), .C2 (n_6_1_553));
INV_X1 i_6_1_33 (.ZN (n_17), .A (n_6_1_16));
AOI222_X1 i_6_1_32 (.ZN (n_6_1_15), .A1 (n_6_959), .A2 (slo___n23232), .B1 (n_6_991)
    , .B2 (slo___n23218), .C1 (n_6_2448), .C2 (n_6_1_588));
INV_X1 i_6_1_31 (.ZN (n_16), .A (n_6_1_15));
AOI222_X1 i_6_1_30 (.ZN (n_6_1_14), .A1 (n_6_895), .A2 (slo___n23367), .B1 (n_6_927)
    , .B2 (n_6_1_625), .C1 (n_6_2479), .C2 (n_6_1_623));
INV_X1 i_6_1_29 (.ZN (n_15), .A (n_6_1_14));
AOI222_X1 i_6_1_28 (.ZN (n_6_1_13), .A1 (n_6_831), .A2 (slo___n23463), .B1 (n_6_863)
    , .B2 (n_6_1_660), .C1 (n_6_2510), .C2 (n_6_1_658));
INV_X1 i_6_1_27 (.ZN (n_14), .A (n_6_1_13));
AOI222_X1 i_6_1_26 (.ZN (n_6_1_12), .A1 (n_6_767), .A2 (n_6_1_694), .B1 (n_6_799)
    , .B2 (n_6_1_695), .C1 (n_6_2541), .C2 (n_6_1_693));
INV_X1 i_6_1_25 (.ZN (n_13), .A (n_6_1_12));
AOI222_X1 i_6_1_24 (.ZN (n_6_1_11), .A1 (n_6_703), .A2 (n_6_1_729), .B1 (n_6_735)
    , .B2 (n_6_1_730), .C1 (n_6_2572), .C2 (n_6_1_728));
INV_X1 i_6_1_23 (.ZN (n_12), .A (n_6_1_11));
AOI222_X1 i_6_1_22 (.ZN (n_6_1_10), .A1 (n_6_639), .A2 (n_6_1_764), .B1 (n_6_671)
    , .B2 (n_6_1_765), .C1 (CLOCK_slo___n64354), .C2 (n_6_1_763));
INV_X1 i_6_1_21 (.ZN (n_11), .A (n_6_1_10));
AOI222_X1 i_6_1_20 (.ZN (n_6_1_9), .A1 (n_6_575), .A2 (n_6_1_799), .B1 (n_6_607), .B2 (n_6_1_800)
    , .C1 (n_6_2634), .C2 (n_6_1_798));
INV_X1 i_6_1_19 (.ZN (n_10), .A (n_6_1_9));
AOI222_X1 i_6_1_18 (.ZN (n_6_1_8), .A1 (n_6_511), .A2 (n_6_1_834), .B1 (n_6_543), .B2 (n_6_1_835)
    , .C1 (n_6_2665), .C2 (CLOCK_sgo__n46922));
INV_X1 i_6_1_17 (.ZN (n_9), .A (n_6_1_8));
AOI222_X1 i_6_1_16 (.ZN (n_6_1_7), .A1 (n_6_447), .A2 (n_6_1_869), .B1 (n_6_479), .B2 (n_6_1_870)
    , .C1 (n_6_2696), .C2 (n_6_1_868));
INV_X1 i_6_1_15 (.ZN (n_8), .A (n_6_1_7));
AOI222_X1 i_6_1_14 (.ZN (n_6_1_6), .A1 (n_6_383), .A2 (n_6_1_904), .B1 (n_6_415), .B2 (n_6_1_905)
    , .C1 (n_6_2727), .C2 (CLOCK_sgo__n46934));
INV_X1 i_6_1_13 (.ZN (n_7), .A (n_6_1_6));
AOI222_X1 i_6_1_12 (.ZN (n_6_1_5), .A1 (n_6_319), .A2 (n_6_1_939), .B1 (n_6_351), .B2 (n_6_1_940)
    , .C1 (n_6_2758), .C2 (CLOCK_sgo__n46937));
INV_X1 i_6_1_11 (.ZN (n_6), .A (n_6_1_5));
AOI222_X1 i_6_1_10 (.ZN (n_6_1_4), .A1 (n_6_255), .A2 (n_6_1_974), .B1 (n_6_287), .B2 (n_6_1_975)
    , .C1 (n_6_2789), .C2 (n_6_1_973));
INV_X1 i_6_1_9 (.ZN (n_5), .A (n_6_1_4));
AOI222_X1 i_6_1_8 (.ZN (n_6_1_3), .A1 (n_6_191), .A2 (n_6_1_1009), .B1 (n_6_223), .B2 (n_6_1_1010)
    , .C1 (n_6_2820), .C2 (CLOCK_sgo__n46950));
INV_X1 i_6_1_7 (.ZN (n_4), .A (n_6_1_3));
AOI222_X1 i_6_1_6 (.ZN (n_6_1_2), .A1 (n_6_127), .A2 (n_6_1_1044), .B1 (n_6_159), .B2 (n_6_1_1045)
    , .C1 (n_6_2851), .C2 (CLOCK_sgo__n46945));
INV_X1 i_6_1_5 (.ZN (n_3), .A (n_6_1_2));
AOI222_X1 i_6_1_4 (.ZN (n_6_1_1), .A1 (n_6_63), .A2 (n_6_1_1079), .B1 (n_6_95), .B2 (n_6_1_1080)
    , .C1 (CLOCK_spw__n65836), .C2 (slo__n13799));
INV_X1 i_6_1_3 (.ZN (n_2), .A (n_6_1_1));
AOI222_X1 i_6_1_2 (.ZN (n_6_1_0), .A1 (slo__n31700), .A2 (opt_ipo_n24358), .B1 (sgo__n1276)
    , .B2 (slo__n30589), .C1 (n_6_31), .C2 (n_6_1_1114));
INV_X1 i_6_1_1 (.ZN (n_1), .A (n_6_1_0));
AND2_X1 i_6_1_0 (.ZN (n_0), .A1 (Multiplicand[0]), .A2 (sgo__n1276));
datapath__0_247 i_6_123 (.p_2 ({n_6_1982, n_6_1981, n_6_1980, n_6_1979, n_6_1978, 
    n_6_1977, n_6_1976, n_6_1975, n_6_1974, n_6_1973, n_6_1972, n_6_1971, n_6_1970, 
    n_6_1969, n_6_1968, n_6_1967, n_6_1966, n_6_1965, n_6_1964, n_6_1963, n_6_1962, 
    n_6_1961, n_6_1960, n_6_1959, n_6_1958, n_6_1957, n_6_1956, n_6_1955, n_6_1954, 
    n_6_1953, n_6_1952, n_6_1951}), .p_0 ({n_6_30, hfn_ipo_n30, drc_ipo_n26573, drc_ipo_n26574, 
    n_6_26, n_6_25, n_6_24, n_6_23, drc_ipo_n26576, drc_ipo_n26577, drc_ipo_n26579, 
    drc_ipo_n26581, drc_ipo_n26582, drc_ipo_n26583, drc_ipo_n26585, drc_ipo_n26584, 
    drc_ipo_n26586, drc_ipo_n26587, drc_ipo_n26588, drc_ipo_n26589, drc_ipo_n26592, 
    drc_ipo_n26590, n_6_8, slo__n4932, n_6_6, slo__n3834, slo__n16572, slo__n3796, 
    slo__n3800, slo__n16608, slo__n5306, sgo__n1276}), .p_1 ({uc_60, n_6_2013, n_6_2012, 
    n_6_2011, n_6_2010, n_6_2009, slo__n27410, n_6_2007, CLOCK_slo__n57743, slo__n40097, 
    n_6_2004, n_6_2003, n_6_2002, n_6_2001, n_6_2000, n_6_1999, n_6_1998, n_6_1997, 
    n_6_1996, n_6_1995, n_6_1994, spw__n68268, CLOCK_slo__n58099, n_6_1_74, n_6_1990, 
    n_6_1989, n_6_1988, slo__n10734, n_6_1986, n_6_1985, n_6_1984, n_6_1983}), .p_1_25_PP_0 (slo__n27410)
    , .p_1_25_PP_1 (slo__n27411));
datapath__0_246 i_6_122 (.p_1 ({n_6_1950, n_6_1949, n_6_1948, n_6_1947, n_6_1946, 
    n_6_1945, n_6_1944, n_6_1943, n_6_1942, n_6_1941, n_6_1940, n_6_1939, n_6_1938, 
    n_6_1937, n_6_1936, n_6_1935, n_6_1934, n_6_1933, n_6_1932, n_6_1931, n_6_1930, 
    n_6_1929, n_6_1928, n_6_1927, n_6_1926, n_6_1925, n_6_1924, n_6_1923, n_6_1922, 
    n_6_1921, n_6_1920, n_6_1919}), .Multiplier ({Multiplier[31], hfn_ipo_n25, drc_ipo_n26625, 
    Multiplier[28], drc_ipoPP_7, Multiplier[26], Multiplier[25], Multiplier[24], 
    drc_ipo_n26618, Multiplier[22], drc_ipo_n26616, Multiplier[20], drc_ipo_n26614, 
    drc_ipo_n26613, Multiplier[17], Multiplier[16], drc_ipo_n26610, Multiplier[14], 
    Multiplier[13], drc_ipo_n26607, drc_ipo_n26606, Multiplier[10], Multiplier[9], 
    Multiplier[8], Multiplier[7], slo__n11938, slo__n4958, slo__n4944, slo__n3804, 
    sgo__n1306, slo__n18930, sgo__n1276}), .p_0 ({uc_59, slo__n40090, n_6_2012, n_6_2011, 
    n_6_2010, n_6_2009, slo__n27410, n_6_2007, n_6_2006, slo__n40097, n_6_2004, n_6_2003, 
    n_6_2002, n_6_2001, n_6_2000, n_6_1999, n_6_1998, n_6_1997, n_6_1996, n_6_1995, 
    n_6_1994, n_6_1993, n_6_1992, n_6_1_74, n_6_1990, n_6_1989, n_6_1988, n_6_1987, 
    slo__n13290, n_6_1985, n_6_1984, n_6_1983}), .drc_ipoPP_0 (drc_ipo_n26624));
datapath__0_242 i_6_119 (.p_2 ({n_6_1918, n_6_1917, n_6_1916, n_6_1915, n_6_1914, 
    n_6_1913, n_6_1912, n_6_1911, n_6_1910, n_6_1909, n_6_1908, n_6_1907, n_6_1906, 
    n_6_1905, n_6_1904, n_6_1903, n_6_1902, n_6_1901, n_6_1900, n_6_1899, n_6_1898, 
    n_6_1897, n_6_1896, n_6_1895, n_6_1894, n_6_1893, n_6_1892, n_6_1891, n_6_1890, 
    n_6_1889, n_6_1888, n_6_1887}), .p_0 ({n_6_30, hfn_ipo_n30, drc_ipo_n26573, drc_ipo_n26574, 
    n_6_26, n_6_25, n_6_24, n_6_23, drc_ipo_n26576, drc_ipo_n26577, drc_ipo_n26579, 
    drc_ipo_n26581, drc_ipo_n26582, drc_ipo_n26583, drc_ipo_n26585, drc_ipo_n26584, 
    drc_ipo_n26586, drc_ipo_n26587, drc_ipo_n26588, drc_ipo_n26589, drc_ipo_n26592, 
    drc_ipo_n26590, n_6_8, slo__n4932, n_6_6, slo__n3834, slo__n16572, slo__n3796, 
    slo__n3800, slo__n16608, slo__n5306, sgo__n1276}), .p_1 ({uc_58, n_6_2044, n_6_2043, 
    n_6_2042, CLOCK_slo__n57242, n_6_2040, slo__n15969, opt_ipo_n45107, slo__n17713, 
    slo__n17680, slo__n17921, slo__n15879, slo__n14104, slo__n39345, n_6_2031, slo___n15411, 
    slo__n28070, CLOCK_opt_ipo_n45744, n_6_2027, n_6_2026, n_6_2025, n_6_2024, n_6_2023, 
    n_6_2022, n_6_2021, opt_ipo_n24075, n_6_2019, n_6_2018, n_6_2017, n_6_2016, n_6_2015, 
    n_6_2014}), .opt_ipoPP_1 (opt_ipo_n24196), .opt_ipoPP_11 (n_6_2021));
datapath__0_241 i_6_118 (.p_1 ({n_6_1886, n_6_1885, n_6_1884, n_6_1883, n_6_1882, 
    n_6_1881, n_6_1880, n_6_1879, n_6_1878, n_6_1877, n_6_1876, n_6_1875, n_6_1874, 
    n_6_1873, n_6_1872, n_6_1871, n_6_1870, n_6_1869, n_6_1868, n_6_1867, n_6_1866, 
    n_6_1865, n_6_1864, n_6_1863, n_6_1862, n_6_1861, n_6_1860, n_6_1859, n_6_1858, 
    n_6_1857, n_6_1856, n_6_1855}), .Multiplier ({Multiplier[31], hfn_ipo_n25, drc_ipo_n26625, 
    drc_ipo_n26624, drc_ipoPP_7, Multiplier[26], Multiplier[25], Multiplier[24], 
    drc_ipo_n26618, Multiplier[22], drc_ipo_n26616, Multiplier[20], drc_ipo_n26614, 
    drc_ipo_n26613, Multiplier[17], Multiplier[16], drc_ipo_n26610, Multiplier[14], 
    Multiplier[13], drc_ipo_n26607, drc_ipo_n26606, Multiplier[10], Multiplier[9], 
    Multiplier[8], Multiplier[7], slo__n11938, slo__n4958, slo__n4944, slo__n3804, 
    sgo__n1306, slo__n18930, sgo__n1276}), .p_0 ({uc_57, n_6_2044, n_6_2043, slo__n39745, 
    n_6_2041, slo__n16063, n_6_2039, opt_ipo_n45107, n_6_2037, n_6_2036, n_6_2035, 
    n_6_2034, n_6_2033, n_6_2032, n_6_2031, slo___n15411, slo__n28070, CLOCK_opt_ipo_n45742, 
    opt_ipo_n24196, n_6_2026, n_6_2025, n_6_2024, n_6_2023, n_6_2022, n_6_2021, opt_ipo_n24075, 
    n_6_2019, n_6_2018, n_6_2017, n_6_2016, n_6_2015, n_6_2014}), .p_0_16_PP_0 (slo___n15411)
    , .p_0_16_PP_1 (slo___n15411), .p_0_15_PP_0 (slo__n28070));
datapath__0_237 i_6_115 (.p_2 ({n_6_1854, n_6_1853, n_6_1852, n_6_1851, n_6_1850, 
    n_6_1849, n_6_1848, n_6_1847, n_6_1846, n_6_1845, n_6_1844, n_6_1843, n_6_1842, 
    n_6_1841, n_6_1840, n_6_1839, n_6_1838, n_6_1837, n_6_1836, n_6_1835, n_6_1834, 
    n_6_1833, n_6_1832, n_6_1831, n_6_1830, n_6_1829, n_6_1828, n_6_1827, n_6_1826, 
    n_6_1825, n_6_1824, n_6_1823}), .p_0 ({n_6_30, hfn_ipo_n30, drc_ipo_n26573, drc_ipo_n26574, 
    n_6_26, n_6_25, n_6_24, n_6_23, drc_ipo_n26576, drc_ipo_n26577, drc_ipo_n26579, 
    drc_ipo_n26581, drc_ipo_n26582, drc_ipo_n26583, drc_ipo_n26585, drc_ipo_n26584, 
    drc_ipo_n26586, drc_ipo_n26587, drc_ipo_n26588, drc_ipo_n26589, drc_ipo_n26592, 
    drc_ipo_n26590, n_6_8, slo__n4932, n_6_6, slo__n3834, slo__n16572, slo__n3796, 
    slo__n3800, slo__n16608, slo__n5306, sgo__n1276}), .p_1 ({uc_56, n_6_2075, n_6_2074, 
    n_6_2073, n_6_2072, slo__n15870, CLOCK_slo__xsl_n57029, n_6_2069, n_6_2068, n_6_2067, 
    n_6_2066, n_6_2065, n_6_2064, slo__n39284, n_6_2062, n_6_2061, n_6_2060, n_6_1_150, 
    n_6_2058, slo__n15402, slo__n39719, n_6_2055, n_6_2054, n_6_2053, n_6_2052, n_6_2051, 
    n_6_2050, n_6_2049, n_6_2048, n_6_2047, n_6_2046, n_6_2045}));
datapath__0_236 i_6_114 (.p_1 ({n_6_1822, n_6_1821, n_6_1820, n_6_1819, n_6_1818, 
    n_6_1817, n_6_1816, n_6_1815, n_6_1814, n_6_1813, n_6_1812, n_6_1811, n_6_1810, 
    n_6_1809, n_6_1808, n_6_1807, n_6_1806, n_6_1805, n_6_1804, n_6_1803, n_6_1802, 
    n_6_1801, n_6_1800, n_6_1799, n_6_1798, n_6_1797, n_6_1796, n_6_1795, n_6_1794, 
    n_6_1793, n_6_1792, n_6_1791}), .Multiplier ({Multiplier[31], hfn_ipo_n25, drc_ipo_n26625, 
    drc_ipo_n26624, drc_ipoPP_7, Multiplier[26], Multiplier[25], Multiplier[24], 
    drc_ipo_n26618, Multiplier[22], drc_ipo_n26616, Multiplier[20], drc_ipo_n26614, 
    drc_ipo_n26613, Multiplier[17], Multiplier[16], drc_ipo_n26610, Multiplier[14], 
    Multiplier[13], drc_ipo_n26607, drc_ipo_n26606, Multiplier[10], Multiplier[9], 
    Multiplier[8], Multiplier[7], slo__n11938, slo__n4958, slo__n4944, slo__n3804, 
    sgo__n1306, slo__n18930, sgo__n1276}), .p_0 ({uc_55, n_6_2075, slo__n38840, n_6_2073, 
    n_6_2072, n_6_2071, slo___n13100, slo__n16022, slo__n18982, slo__n17671, n_6_2066, 
    slo__n15443, slo__n14771, slo__n39285, slo__n14766, slo__n15745, slo__n36350, 
    n_6_1_150, n_6_2058, n_6_2057, n_6_2056, n_6_2055, n_6_2054, slo__n16524, slo__n15821, 
    n_6_2051, n_6_2050, n_6_2049, slo__n10634, n_6_2047, n_6_2046, n_6_2045}), .p_0_25_PP_0 (slo___n13099));
datapath__0_232 i_6_111 (.p_2 ({n_6_1790, n_6_1789, n_6_1788, n_6_1787, n_6_1786, 
    n_6_1785, n_6_1784, n_6_1783, n_6_1782, n_6_1781, n_6_1780, n_6_1779, n_6_1778, 
    n_6_1777, n_6_1776, n_6_1775, n_6_1774, n_6_1773, n_6_1772, n_6_1771, n_6_1770, 
    n_6_1769, n_6_1768, n_6_1767, n_6_1766, n_6_1765, n_6_1764, n_6_1763, n_6_1762, 
    n_6_1761, n_6_1760, n_6_1759}), .p_0 ({n_6_30, hfn_ipo_n31, drc_ipo_n26573, n_6_27, 
    n_6_26, n_6_25, n_6_24, n_6_23, drc_ipo_n26576, drc_ipo_n26577, drc_ipo_n26579, 
    drc_ipo_n26581, drc_ipo_n26582, drc_ipo_n26583, drc_ipo_n26585, drc_ipo_n26584, 
    drc_ipo_n26586, drc_ipo_n26587, drc_ipo_n26588, drc_ipo_n26589, drc_ipo_n26592, 
    drc_ipo_n26590, n_6_8, slo__n4932, n_6_6, slo__n3834, slo__n16572, slo__n3796, 
    slo__n3800, slo__n16608, slo__n5306, sgo__n1276}), .p_1 ({uc_54, CLOCK_slo__n54289, 
    n_6_2105, slo__n33292, n_6_2103, n_6_2102, n_6_2101, n_6_2100, CLOCK_slo__n56418, 
    n_6_2098, spw__n69101, slo___n13213, slo__n39714, n_6_2094, n_6_2093, slo__n18122, 
    opt_ipo_n24707, n_6_2090, n_6_2089, n_6_2088, n_6_2087, n_6_2086, n_6_2085, slo__sro_n30921, 
    n_6_2083, n_6_2082, n_6_2081, n_6_2080, n_6_2079, n_6_2078, n_6_2077, n_6_2076}));
datapath__0_231 i_6_110 (.p_1 ({n_6_1758, n_6_1757, n_6_1756, n_6_1755, n_6_1754, 
    n_6_1753, n_6_1752, n_6_1751, n_6_1750, n_6_1749, n_6_1748, n_6_1747, n_6_1746, 
    n_6_1745, n_6_1744, n_6_1743, n_6_1742, n_6_1741, n_6_1740, n_6_1739, n_6_1738, 
    n_6_1737, n_6_1736, n_6_1735, n_6_1734, n_6_1733, n_6_1732, n_6_1731, n_6_1730, 
    n_6_1729, n_6_1728, n_6_1727}), .Multiplier ({Multiplier[31], hfn_ipo_n26, drc_ipo_n26625, 
    drc_ipo_n26624, drc_ipoPP_7, Multiplier[26], Multiplier[25], Multiplier[24], 
    drc_ipo_n26618, Multiplier[22], drc_ipo_n26616, drc_ipo_n26615, drc_ipo_n26614, 
    drc_ipo_n26613, Multiplier[17], Multiplier[16], drc_ipo_n26610, Multiplier[14], 
    Multiplier[13], drc_ipo_n26607, drc_ipo_n26606, Multiplier[10], Multiplier[9], 
    Multiplier[8], Multiplier[7], slo__n11938, slo__n4958, slo__n4944, slo__n3804, 
    sgo__n1306, slo__n18930, sgo__n1276}), .p_0 ({uc_53, n_6_2106, n_6_2105, slo__n33292, 
    n_6_2103, n_6_2102, n_6_2101, n_6_2100, slo___n18137, n_6_2098, spw__n69100, 
    slo___n13213, n_6_2095, n_6_2094, n_6_2093, n_6_2092, opt_ipo_n24707, n_6_2090, 
    n_6_2089, n_6_2088, n_6_2087, n_6_2086, n_6_2085, slo__sro_n30921, n_6_2083, 
    n_6_2082, CLOCK_slo__n55073, n_6_2080, n_6_2079, CLOCK_slo__n57293, n_6_2077, 
    n_6_2076}));
datapath__0_227 i_6_107 (.p_2 ({n_6_1726, n_6_1725, n_6_1724, n_6_1723, n_6_1722, 
    n_6_1721, n_6_1720, n_6_1719, n_6_1718, n_6_1717, n_6_1716, n_6_1715, n_6_1714, 
    n_6_1713, n_6_1712, n_6_1711, n_6_1710, n_6_1709, n_6_1708, n_6_1707, n_6_1706, 
    n_6_1705, n_6_1704, n_6_1703, n_6_1702, n_6_1701, n_6_1700, n_6_1699, n_6_1698, 
    n_6_1697, n_6_1696, n_6_1695}), .p_0 ({n_6_30, hfn_ipo_n31, drc_ipo_n26573, drc_ipo_n26574, 
    n_6_26, n_6_25, n_6_24, n_6_23, drc_ipo_n26576, drc_ipo_n26577, drc_ipo_n26579, 
    drc_ipo_n26581, drc_ipo_n26582, drc_ipo_n26583, drc_ipo_n26585, drc_ipo_n26584, 
    drc_ipo_n26586, drc_ipo_n26587, drc_ipo_n26588, drc_ipo_n26589, drc_ipo_n26592, 
    drc_ipo_n26590, n_6_8, slo__n4932, n_6_6, slo__n3834, slo__n16572, slo__n3796, 
    slo__n3800, slo__n16608, slo__n5306, hfn_ipo_n29}), .p_1 ({uc_52, n_6_2137, n_6_2136, 
    n_6_2135, n_6_2134, n_6_2133, n_6_2132, slo__n30795, slo__n18328, opt_ipo_n45324, 
    n_6_2128, n_6_2127, n_6_2126, n_6_2125, slo__n15420, n_6_2123, n_6_2122, n_6_2121, 
    n_6_2120, n_6_2119, opt_ipo_n24541, n_6_2117, n_6_2116, n_6_2115, n_6_2114, n_6_2113, 
    n_6_2112, n_6_2111, n_6_2110, n_6_2109, n_6_2108, n_6_2107}), .p_1_22_PP_5 (opt_ipo_n45324));
datapath__0_226 i_6_106 (.p_1 ({n_6_1694, n_6_1693, n_6_1692, n_6_1691, n_6_1690, 
    n_6_1689, n_6_1688, n_6_1687, n_6_1686, n_6_1685, n_6_1684, n_6_1683, n_6_1682, 
    n_6_1681, n_6_1680, n_6_1679, n_6_1678, n_6_1677, n_6_1676, n_6_1675, n_6_1674, 
    n_6_1673, n_6_1672, n_6_1671, n_6_1670, n_6_1669, n_6_1668, n_6_1667, n_6_1666, 
    n_6_1665, n_6_1664, n_6_1663}), .Multiplier ({Multiplier[31], hfn_ipo_n26, drc_ipo_n26625, 
    drc_ipo_n26624, drc_ipoPP_7, Multiplier[26], Multiplier[25], Multiplier[24], 
    drc_ipo_n26618, Multiplier[22], drc_ipo_n26616, drc_ipo_n26615, drc_ipo_n26614, 
    drc_ipo_n26613, Multiplier[17], Multiplier[16], drc_ipo_n26610, Multiplier[14], 
    Multiplier[13], drc_ipo_n26607, drc_ipo_n26606, Multiplier[10], Multiplier[9], 
    Multiplier[8], Multiplier[7], slo__n11938, slo__n4958, slo__n4944, slo__n3804, 
    sgo__n1306, slo__n18930, hfn_ipo_n29}), .p_0 ({uc_51, n_6_2137, n_6_2136, n_6_2135, 
    slo__n14143, n_6_2133, n_6_2132, slo__n30795, n_6_2130, opt_ipo_n45324, slo__n13394, 
    n_6_2127, n_6_2126, n_6_2125, n_6_2124, n_6_2123, n_6_2122, n_6_2121, n_6_2120, 
    n_6_2119, opt_ipo_n24541, n_6_2117, n_6_2116, n_6_2115, n_6_2114, n_6_2113, n_6_2112, 
    n_6_2111, n_6_2110, n_6_2109, n_6_2108, n_6_2107}), .p_0_24_PP_1 (slo__n30795));
datapath__0_222 i_6_103 (.p_2 ({n_6_1662, n_6_1661, n_6_1660, n_6_1659, n_6_1658, 
    n_6_1657, n_6_1656, n_6_1655, n_6_1654, n_6_1653, n_6_1652, n_6_1651, n_6_1650, 
    n_6_1649, n_6_1648, n_6_1647, n_6_1646, n_6_1645, n_6_1644, n_6_1643, n_6_1642, 
    n_6_1641, n_6_1640, n_6_1639, n_6_1638, n_6_1637, n_6_1636, n_6_1635, n_6_1634, 
    n_6_1633, n_6_1632, n_6_1631}), .p_0 ({n_6_30, hfn_ipo_n31, drc_ipo_n26573, drc_ipo_n26574, 
    n_6_26, n_6_25, n_6_24, n_6_23, drc_ipo_n26576, drc_ipo_n26577, drc_ipo_n26579, 
    drc_ipo_n26581, drc_ipo_n26582, drc_ipo_n26583, drc_ipo_n26585, drc_ipo_n26584, 
    drc_ipo_n26586, drc_ipo_n26587, drc_ipo_n26588, drc_ipo_n26589, drc_ipo_n26592, 
    drc_ipo_n26590, n_6_8, slo__n4932, slo__n26805, slo__n26713, slo__n16572, slo__n3796, 
    slo__n3800, slo__n16608, slo__n5306, hfn_ipo_n29}), .p_1 ({uc_50, n_6_2168, n_6_2167, 
    n_6_2166, n_6_2165, n_6_2164, n_6_2163, n_6_2162, n_6_2161, n_6_2160, n_6_2159, 
    n_6_2158, n_6_2157, slo___n13169, n_6_2155, n_6_2154, n_6_2153, CLOCK_slo__n54674, 
    n_6_2151, slo__n28104, n_6_2149, n_6_2148, n_6_2147, n_6_2146, n_6_2145, n_6_2144, 
    n_6_2143, n_6_2142, n_6_2141, n_6_2140, n_6_2139, n_6_2138}), .opt_ipoPP_5 (n_6_2158));
datapath__0_221 i_6_102 (.p_1 ({n_6_1630, n_6_1629, n_6_1628, n_6_1627, n_6_1626, 
    n_6_1625, n_6_1624, n_6_1623, n_6_1622, n_6_1621, n_6_1620, n_6_1619, n_6_1618, 
    n_6_1617, n_6_1616, n_6_1615, n_6_1614, n_6_1613, n_6_1612, n_6_1611, n_6_1610, 
    n_6_1609, n_6_1608, n_6_1607, n_6_1606, n_6_1605, n_6_1604, n_6_1603, n_6_1602, 
    n_6_1601, n_6_1600, n_6_1599}), .Multiplier ({Multiplier[31], hfn_ipo_n26, drc_ipo_n26625, 
    drc_ipo_n26624, drc_ipoPP_7, Multiplier[26], Multiplier[25], Multiplier[24], 
    drc_ipo_n26618, Multiplier[22], drc_ipo_n26616, drc_ipo_n26615, drc_ipo_n26614, 
    drc_ipo_n26613, Multiplier[17], Multiplier[16], drc_ipo_n26610, Multiplier[14], 
    CLOCK_sgo__n46814, drc_ipo_n26607, drc_ipo_n26606, Multiplier[10], Multiplier[9], 
    Multiplier[8], Multiplier[7], slo__n11938, slo__n4958, slo__n4944, slo__n3804, 
    sgo__n1306, slo__n18930, hfn_ipo_n29}), .p_0 ({uc_49, n_6_2168, n_6_2167, slo__n15903, 
    slo__n15894, slo__n15930, n_6_2163, n_6_2162, n_6_2161, n_6_2160, n_6_2159, n_6_2158, 
    n_6_2157, slo__n14207, slo__n13153, n_6_2154, n_6_2153, n_6_2152, slo__n19320, 
    slo__n28104, n_6_2149, n_6_2148, n_6_2147, n_6_2146, n_6_2145, n_6_2144, n_6_2143, 
    n_6_2142, n_6_2141, n_6_2140, n_6_2139, n_6_2138}));
datapath__0_217 i_6_99 (.p_2 ({n_6_1598, n_6_1597, n_6_1596, n_6_1595, n_6_1594, 
    n_6_1593, n_6_1592, n_6_1591, n_6_1590, n_6_1589, n_6_1588, n_6_1587, n_6_1586, 
    n_6_1585, n_6_1584, n_6_1583, n_6_1582, n_6_1581, n_6_1580, n_6_1579, n_6_1578, 
    n_6_1577, n_6_1576, n_6_1575, n_6_1574, n_6_1573, n_6_1572, n_6_1571, n_6_1570, 
    n_6_1569, n_6_1568, n_6_1567}), .p_0 ({n_6_30, hfn_ipo_n32, drc_ipo_n26573, drc_ipo_n26574, 
    n_6_26, n_6_25, n_6_24, n_6_23, drc_ipo_n26576, drc_ipo_n26577, drc_ipo_n26579, 
    drc_ipo_n26581, drc_ipo_n26582, drc_ipo_n26583, drc_ipo_n26585, drc_ipo_n26584, 
    drc_ipo_n26586, drc_ipo_n26587, drc_ipo_n26588, drc_ipo_n26589, drc_ipo_n26592, 
    drc_ipo_n26590, slo__n26638, slo__n4932, slo__n26805, slo__n26713, slo__n16572, 
    slo__n3796, slo__n3800, slo__n16608, slo__n31700, hfn_ipo_n29}), .p_1 ({uc_48, 
    n_6_2199, n_6_2198, n_6_2197, n_6_2196, n_6_2195, opt_ipo_n45121, n_6_2193, n_6_2192, 
    n_6_2191, n_6_2190, n_6_2189, slo___n17633, n_6_2187, n_6_2186, n_6_2185, n_6_2184, 
    slo__n38240, n_6_2182, n_6_2181, n_6_2180, n_6_2179, n_6_2178, n_6_2177, n_6_2176, 
    CLOCK_opt_ipo_n45969, n_6_2174, n_6_2173, CLOCK_opt_ipo_n45779, n_6_2171, n_6_2170, 
    n_6_2169}));
datapath__0_216 i_6_98 (.p_1 ({n_6_1566, n_6_1565, n_6_1564, n_6_1563, n_6_1562, 
    n_6_1561, n_6_1560, n_6_1559, n_6_1558, n_6_1557, n_6_1556, n_6_1555, n_6_1554, 
    n_6_1553, n_6_1552, n_6_1551, n_6_1550, n_6_1549, n_6_1548, n_6_1547, n_6_1546, 
    n_6_1545, n_6_1544, n_6_1543, n_6_1542, n_6_1541, n_6_1540, n_6_1539, n_6_1538, 
    n_6_1537, n_6_1536, n_6_1535}), .Multiplier ({Multiplier[31], hfn_ipo_n26, drc_ipo_n26625, 
    drc_ipo_n26624, drc_ipoPP_7, Multiplier[26], Multiplier[25], Multiplier[24], 
    drc_ipo_n26618, Multiplier[22], drc_ipo_n26616, drc_ipo_n26615, drc_ipo_n26614, 
    drc_ipo_n26613, Multiplier[17], Multiplier[16], drc_ipo_n26610, drc_ipo_n26609, 
    CLOCK_sgo__n46814, drc_ipo_n26607, drc_ipo_n26606, Multiplier[10], Multiplier[9], 
    Multiplier[8], Multiplier[7], slo__n11938, slo__n4958, slo__n4944, slo__n3804, 
    sgo__n1306, slo__n18930, hfn_ipo_n29}), .p_0 ({uc_47, n_6_2199, n_6_2198, slo__n14019, 
    n_6_2196, n_6_2195, opt_ipo_n45121, CLOCK_slo__n57308, n_6_2192, n_6_2191, n_6_2190, 
    n_6_2189, slo__n11671, slo__n12943, n_6_2186, n_6_2185, n_6_2184, n_6_2183, n_6_2182, 
    n_6_2181, slo__n39452, n_6_2179, n_6_2178, n_6_2177, n_6_2176, CLOCK_opt_ipo_n45969, 
    n_6_2174, n_6_2173, CLOCK_opt_ipo_n45779, n_6_2171, n_6_2170, n_6_2169}), .Multiplier_13_PP_0 (CLOCK_sgo__n46814));
datapath__0_212 i_6_95 (.p_2 ({n_6_1534, n_6_1533, n_6_1532, n_6_1531, n_6_1530, 
    n_6_1529, n_6_1528, n_6_1527, n_6_1526, n_6_1525, n_6_1524, n_6_1523, n_6_1522, 
    n_6_1521, n_6_1520, n_6_1519, n_6_1518, n_6_1517, n_6_1516, n_6_1515, n_6_1514, 
    n_6_1513, n_6_1512, n_6_1511, n_6_1510, n_6_1509, n_6_1508, n_6_1507, n_6_1506, 
    n_6_1505, n_6_1504, n_6_1503}), .p_0 ({n_6_30, hfn_ipo_n32, drc_ipo_n26573, drc_ipo_n26574, 
    n_6_26, n_6_25, n_6_24, n_6_23, drc_ipo_n26576, drc_ipo_n26577, drc_ipo_n26579, 
    drc_ipo_n26581, drc_ipo_n26582, drc_ipo_n26583, drc_ipo_n26585, drc_ipo_n26584, 
    drc_ipo_n26586, drc_ipo_n26587, drc_ipo_n26588, drc_ipo_n26589, drc_ipo_n26592, 
    drc_ipo_n26590, slo__n26638, slo__n4932, slo__n26805, slo__n26713, slo__n16572, 
    slo__n26761, slo__n3800, slo__n16608, slo__n31700, hfn_ipo_n29}), .p_1 ({uc_46, 
    n_6_2230, n_6_2229, n_6_2228, slo___n15724, slo__sro_n2968, n_6_2225, n_6_2224, 
    n_6_2223, n_6_2222, n_6_2221, n_6_2220, n_6_2219, opt_ipo_n24721, n_6_2217, n_6_2216, 
    n_6_2215, slo__n12843, slo__n14640, n_6_2212, n_6_2211, n_6_2210, n_6_2209, n_6_2208, 
    n_6_2207, n_6_2206, n_6_2205, n_6_2204, n_6_2203, n_6_2202, CLOCK_opt_ipo_n45894, 
    n_6_2200}), .opt_ipoPP_2 (CLOCK_opt_ipo_n45893));
datapath__0_211 i_6_94 (.p_1 ({n_6_1502, n_6_1501, n_6_1500, n_6_1499, n_6_1498, 
    n_6_1497, n_6_1496, n_6_1495, n_6_1494, n_6_1493, n_6_1492, n_6_1491, n_6_1490, 
    n_6_1489, n_6_1488, n_6_1487, n_6_1486, n_6_1485, n_6_1484, n_6_1483, n_6_1482, 
    n_6_1481, n_6_1480, n_6_1479, n_6_1478, n_6_1477, n_6_1476, n_6_1475, n_6_1474, 
    n_6_1473, n_6_1472, n_6_1471}), .Multiplier ({Multiplier[31], hfn_ipo_n27, drc_ipo_n26625, 
    drc_ipo_n26624, drc_ipoPP_7, Multiplier[26], Multiplier[25], Multiplier[24], 
    drc_ipo_n26618, drc_ipo_n26617, drc_ipo_n26616, drc_ipo_n26615, drc_ipo_n26614, 
    drc_ipo_n26613, Multiplier[17], Multiplier[16], drc_ipo_n26610, drc_ipo_n26609, 
    CLOCK_sgo__n46814, drc_ipo_n26607, drc_ipo_n26606, Multiplier[10], Multiplier[9], 
    Multiplier[8], Multiplier[7], slo__n11938, slo__n4958, slo__n4944, slo__n3804, 
    sgo__n1306, slo__n18930, hfn_ipo_n29}), .p_0 ({uc_45, n_6_2230, n_6_2229, n_6_2228, 
    slo__n14647, slo__sro_n2968, n_6_2225, n_6_2224, CLOCK_slo__n53754, n_6_2222, 
    n_6_2221, n_6_2220, slo__n39406, CLOCK_slo__n53479, slo__n38973, n_6_2216, slo__n16143, 
    n_6_2214, n_6_2213, n_6_2212, n_6_2211, n_6_2210, n_6_2209, n_6_2208, n_6_2207, 
    n_6_2206, n_6_2205, n_6_2204, n_6_2203, n_6_2202, CLOCK_opt_ipo_n45893, n_6_2200})
    , .drc_ipoPP_0 (drc_ipo_n26602));
datapath__0_207 i_6_91 (.p_2 ({n_6_1470, n_6_1469, n_6_1468, n_6_1467, n_6_1466, 
    n_6_1465, n_6_1464, n_6_1463, n_6_1462, n_6_1461, n_6_1460, n_6_1459, n_6_1458, 
    n_6_1457, n_6_1456, n_6_1455, n_6_1454, n_6_1453, n_6_1452, n_6_1451, n_6_1450, 
    n_6_1449, n_6_1448, n_6_1447, n_6_1446, n_6_1445, n_6_1444, n_6_1443, n_6_1442, 
    n_6_1441, n_6_1440, n_6_1439}), .p_0 ({n_6_30, hfn_ipo_n32, drc_ipo_n26573, drc_ipo_n26574, 
    n_6_26, n_6_25, drc_ipo_n26575, CLOCK_sgo__n47049, drc_ipo_n26576, drc_ipo_n26577, 
    drc_ipo_n26579, drc_ipo_n26581, drc_ipo_n26582, drc_ipo_n26583, drc_ipo_n26585, 
    drc_ipo_n26584, drc_ipo_n26586, drc_ipo_n26587, drc_ipo_n26588, drc_ipo_n26589, 
    drc_ipo_n26592, drc_ipo_n26590, slo__n26638, slo__n4932, slo__n26805, slo__n26713, 
    slo__n16572, slo__n26761, slo__n3800, slo__n16608, slo__n31700, hfn_ipo_n29})
    , .p_1 ({uc_44, n_6_2261, n_6_2260, n_6_2259, n_6_2258, n_6_2257, n_6_2256, n_6_2255, 
    slo__n17378, n_6_2253, n_6_2252, opt_ipo_n24431, n_6_2250, n_6_2249, n_6_2248, 
    n_6_2247, n_6_2246, n_6_2245, n_6_2244, n_6_2243, n_6_2242, n_6_2241, n_6_2240, 
    CLOCK_opt_ipo_n45978, n_6_2238, n_6_2237, n_6_2236, n_6_2235, n_6_2234, n_6_2233, 
    CLOCK_slo__n55465, n_6_2231}));
datapath__0_206 i_6_90 (.p_1 ({n_6_1438, n_6_1437, n_6_1436, n_6_1435, n_6_1434, 
    n_6_1433, n_6_1432, n_6_1431, n_6_1430, n_6_1429, n_6_1428, n_6_1427, n_6_1426, 
    n_6_1425, n_6_1424, n_6_1423, n_6_1422, n_6_1421, n_6_1420, n_6_1419, n_6_1418, 
    n_6_1417, n_6_1416, n_6_1415, n_6_1414, n_6_1413, n_6_1412, n_6_1411, n_6_1410, 
    n_6_1409, n_6_1408, n_6_1407}), .Multiplier ({Multiplier[31], hfn_ipo_n27, drc_ipo_n26625, 
    drc_ipo_n26624, drc_ipoPP_7, Multiplier[26], drc_ipo_n26621, drc_ipo_n26620, 
    drc_ipo_n26618, drc_ipo_n26617, drc_ipo_n26616, drc_ipo_n26615, drc_ipo_n26614, 
    drc_ipo_n26613, drc_ipoPP_4, Multiplier[16], drc_ipo_n26610, drc_ipo_n26609, 
    CLOCK_sgo__n46814, drc_ipo_n26607, drc_ipo_n26606, Multiplier[10], drc_ipoPP_1, 
    Multiplier[8], drc_ipo_n26602, slo__n11938, drc_ipo_n26600, slo__n4944, slo__n3804, 
    sgo__n1306, slo__n18930, hfn_ipo_n29}), .p_0 ({uc_43, n_6_2261, n_6_2260, n_6_2259, 
    slo__n18019, n_6_2257, slo__n17416, n_6_2255, n_6_2254, n_6_2253, n_6_2252, opt_ipo_n24431, 
    n_6_2250, n_6_2249, n_6_2248, slo__n39417, slo__n11990, slo__n14684, slo__n16747, 
    n_6_2243, n_6_2242, n_6_2241, slo__n14568, CLOCK_opt_ipo_n45978, n_6_2238, n_6_2237, 
    slo__n17088, CLOCK_slo__n58195, n_6_2234, n_6_2233, n_6_2232, n_6_2231}), .drc_ipoPP_0 (drc_ipo_n26599)
    , .drc_ipoPP_1 (drc_ipoPP_0), .drc_ipoPP_2 (CLOCK_sgo__n46808));
datapath__0_202 i_6_87 (.p_2 ({n_6_1406, n_6_1405, n_6_1404, n_6_1403, n_6_1402, 
    n_6_1401, n_6_1400, n_6_1399, n_6_1398, n_6_1397, n_6_1396, n_6_1395, n_6_1394, 
    n_6_1393, n_6_1392, n_6_1391, n_6_1390, n_6_1389, n_6_1388, n_6_1387, n_6_1386, 
    n_6_1385, n_6_1384, n_6_1383, n_6_1382, n_6_1381, n_6_1380, n_6_1379, n_6_1378, 
    n_6_1377, n_6_1376, n_6_1375}), .p_0 ({n_6_30, hfn_ipo_n32, drc_ipo_n26573, drc_ipo_n26574, 
    n_6_26, n_6_25, drc_ipo_n26575, CLOCK_sgo__n47049, drc_ipo_n26576, drc_ipo_n26577, 
    drc_ipo_n26579, drc_ipo_n26581, drc_ipo_n26582, drc_ipo_n26583, drc_ipo_n26585, 
    drc_ipo_n26584, drc_ipo_n26586, drc_ipo_n26587, drc_ipo_n26588, drc_ipo_n26589, 
    drc_ipo_n26592, drc_ipo_n26590, slo__n26638, slo__n4932, slo__n26805, slo__n26713, 
    slo__n16572, slo__n26761, slo__n3800, slo__n16608, slo__n31700, hfn_ipo_n29})
    , .p_1 ({uc_42, n_6_2292, n_6_2291, opt_ipo_n24063, n_6_2289, CLOCK_slo__n55658, 
    n_6_2287, n_6_2286, n_6_2285, n_6_2284, n_6_2283, opt_ipo_n24727, n_6_2281, n_6_2280, 
    slo__n32747, n_6_2278, n_6_2277, spw__n67799, n_6_2275, n_6_2274, n_6_2273, slo__n28538, 
    n_6_2271, n_6_2270, n_6_2269, n_6_2268, n_6_2267, n_6_2266, CLOCK_opt_ipo_n45906, 
    CLOCK_opt_ipo_n45803, n_6_2263, n_6_2262}));
datapath__0_201 i_6_86 (.p_1 ({n_6_1374, n_6_1373, n_6_1372, n_6_1371, n_6_1370, 
    n_6_1369, n_6_1368, n_6_1367, n_6_1366, n_6_1365, n_6_1364, n_6_1363, n_6_1362, 
    n_6_1361, n_6_1360, n_6_1359, n_6_1358, n_6_1357, n_6_1356, n_6_1355, n_6_1354, 
    n_6_1353, n_6_1352, n_6_1351, n_6_1350, n_6_1349, n_6_1348, n_6_1347, n_6_1346, 
    n_6_1345, n_6_1344, n_6_1343}), .Multiplier ({Multiplier[31], hfn_ipo_n27, drc_ipo_n26625, 
    drc_ipo_n26624, drc_ipoPP_7, Multiplier[26], drc_ipo_n26621, drc_ipo_n26620, 
    drc_ipo_n26618, drc_ipo_n26617, drc_ipo_n26616, drc_ipo_n26615, drc_ipo_n26614, 
    drc_ipo_n26613, drc_ipoPP_4, CLOCK_sgo__n46808, drc_ipo_n26610, drc_ipo_n26609, 
    CLOCK_sgo__n46814, drc_ipo_n26607, drc_ipo_n26606, Multiplier[10], drc_ipoPP_1, 
    drc_ipoPP_0, drc_ipo_n26602, drc_ipo_n26599, drc_ipo_n26600, slo__n4944, slo__n3804, 
    sgo__n1306, slo__n18930, hfn_ipo_n29}), .p_0 ({uc_41, n_6_2292, n_6_2291, opt_ipo_n24063, 
    n_6_2289, slo___n13086, n_6_2287, n_6_2286, slo__n38193, n_6_2284, CLOCK_slo__n57977, 
    opt_ipo_n24727, slo__n37502, n_6_2280, slo__n32747, n_6_2278, slo__n16450, slo__n18848, 
    slo__n11487, CLOCK_slo__n54187, n_6_2273, slo__n28538, slo__n13303, slo__n17020, 
    slo__n14095, slo__n10929, n_6_2267, n_6_2266, CLOCK_opt_ipo_n45906, CLOCK_opt_ipo_n45803, 
    n_6_2263, n_6_2262}), .p_0_17_PP_1 (slo__n32747), .opt_ipoPP_0 (n_6_2266), .p_0_16_PP_5 (n_6_2278));
datapath__0_197 i_6_83 (.p_2 ({n_6_1342, n_6_1341, n_6_1340, n_6_1339, n_6_1338, 
    n_6_1337, n_6_1336, n_6_1335, n_6_1334, n_6_1333, n_6_1332, n_6_1331, n_6_1330, 
    n_6_1329, n_6_1328, n_6_1327, n_6_1326, n_6_1325, n_6_1324, n_6_1323, n_6_1322, 
    n_6_1321, n_6_1320, n_6_1319, n_6_1318, n_6_1317, n_6_1316, n_6_1315, n_6_1314, 
    n_6_1313, n_6_1312, n_6_1311}), .p_0 ({n_6_30, hfn_ipo_n32, drc_ipo_n26573, drc_ipo_n26574, 
    n_6_26, n_6_25, drc_ipo_n26575, CLOCK_sgo__n47049, drc_ipo_n26576, drc_ipo_n26577, 
    drc_ipo_n26579, drc_ipo_n26581, drc_ipo_n26582, drc_ipo_n26583, drc_ipo_n26585, 
    drc_ipo_n26584, drc_ipo_n26586, drc_ipo_n26587, drc_ipo_n26588, drc_ipo_n26589, 
    drc_ipo_n26592, drc_ipo_n26590, slo__n26638, slo__n4932, slo__n26805, slo__n26713, 
    slo__n16572, slo__n26761, slo__n3800, slo__n16608, slo__n31700, hfn_ipo_n29})
    , .p_1 ({uc_40, n_6_2323, n_6_2322, opt_ipo_n45134, n_6_2320, n_6_2319, n_6_2318, 
    n_6_2317, CLOCK_slo__n57799, n_6_2315, n_6_2314, CLOCK_slo__n54661, slo__n36345, 
    n_6_2311, n_6_2310, n_6_2309, n_6_2308, n_6_2307, n_6_2306, n_6_2305, n_6_2304, 
    n_6_2303, n_6_2302, n_6_2301, slo__n19067, n_6_2299, n_6_2298, n_6_2297, CLOCK_opt_ipo_n45807, 
    n_6_2295, n_6_2294, n_6_2293}), .opt_ipoPP_1 (opt_ipo_n45132));
datapath__0_196 i_6_82 (.p_1 ({n_6_1310, n_6_1309, n_6_1308, n_6_1307, n_6_1306, 
    n_6_1305, n_6_1304, n_6_1303, n_6_1302, n_6_1301, n_6_1300, n_6_1299, n_6_1298, 
    n_6_1297, n_6_1296, n_6_1295, n_6_1294, n_6_1293, n_6_1292, n_6_1291, n_6_1290, 
    n_6_1289, n_6_1288, n_6_1287, n_6_1286, n_6_1285, n_6_1284, n_6_1283, n_6_1282, 
    n_6_1281, n_6_1280, n_6_1279}), .Multiplier ({Multiplier[31], hfn_ipo_n27, drc_ipo_n26625, 
    drc_ipo_n26624, drc_ipoPP_7, Multiplier[26], drc_ipo_n26621, drc_ipo_n26620, 
    drc_ipo_n26618, drc_ipo_n26617, drc_ipo_n26616, drc_ipo_n26615, drc_ipo_n26614, 
    drc_ipo_n26613, drc_ipoPP_4, CLOCK_sgo__n46808, drc_ipo_n26610, drc_ipo_n26609, 
    CLOCK_sgo__n46814, drc_ipo_n26607, drc_ipo_n26606, drc_ipo_n26605, drc_ipoPP_1, 
    drc_ipoPP_0, drc_ipo_n26602, drc_ipo_n26599, drc_ipo_n26600, slo__n4944, slo__n3804, 
    sgo__n1306, drc_ipo_n26598, hfn_ipo_n29}), .p_0 ({uc_39, n_6_2323, n_6_2322, 
    opt_ipo_n45134, CLOCK_slo__n57760, n_6_2319, n_6_2318, n_6_2317, n_6_2316, slo__n37528, 
    n_6_2314, n_6_2313, n_6_2312, n_6_2311, CLOCK_slo__n54206, slo__n18991, n_6_2308, 
    slo__n12014, n_6_2306, n_6_2305, n_6_2304, slo__n17821, n_6_2302, slo__n16529, 
    n_6_2300, n_6_2299, slo__n16348, slo__n11253, CLOCK_slo__n64621, n_6_2295, n_6_2294, 
    n_6_2293}), .opt_ipoPP_1 (n_6_2302));
datapath__0_192 i_6_79 (.p_2 ({n_6_1278, n_6_1277, n_6_1276, n_6_1275, n_6_1274, 
    n_6_1273, n_6_1272, n_6_1271, n_6_1270, n_6_1269, n_6_1268, n_6_1267, n_6_1266, 
    n_6_1265, n_6_1264, n_6_1263, n_6_1262, n_6_1261, n_6_1260, n_6_1259, n_6_1258, 
    n_6_1257, n_6_1256, n_6_1255, n_6_1254, n_6_1253, n_6_1252, n_6_1251, n_6_1250, 
    n_6_1249, n_6_1248, n_6_1247}), .p_0 ({n_6_30, hfn_ipo_n32, drc_ipo_n26573, drc_ipo_n26574, 
    n_6_26, n_6_25, drc_ipo_n26575, CLOCK_sgo__n47049, drc_ipo_n26576, drc_ipo_n26577, 
    drc_ipo_n26579, drc_ipo_n26581, drc_ipo_n26582, drc_ipo_n26583, drc_ipo_n26585, 
    drc_ipo_n26584, drc_ipo_n26586, drc_ipo_n26587, drc_ipo_n26588, drc_ipo_n26589, 
    drc_ipo_n26592, drc_ipo_n26590, slo__n26638, slo__n4932, slo__n26805, slo__n26713, 
    slo__n16572, slo__n26761, slo__n3800, slo__n16608, slo__n31700, hfn_ipo_n29})
    , .p_1 ({uc_38, n_6_2354, opt_ipo_n45138, n_6_2352, n_6_2351, n_6_2350, CLOCK_slo__n55312, 
    slo__n17435, opt_ipo_n43935, n_6_2346, n_6_2345, n_6_2344, n_6_2343, n_6_2342, 
    n_6_2341, n_6_2340, slo__n14603, n_6_2338, n_6_2337, n_6_2336, n_6_2335, n_6_2334, 
    n_6_2333, slo__n13528, opt_ipo_n23778, n_6_2330, n_6_2329, opt_ipo_n26244, slo__n17619, 
    slo__n13728, CLOCK_opt_ipo_n45918, n_6_2324}), .opt_ipoPP_0 (CLOCK_opt_ipo_n46265));
datapath__0_191 i_6_78 (.p_1 ({n_6_1246, n_6_1245, n_6_1244, n_6_1243, n_6_1242, 
    n_6_1241, n_6_1240, n_6_1239, n_6_1238, n_6_1237, n_6_1236, n_6_1235, n_6_1234, 
    n_6_1233, n_6_1232, n_6_1231, n_6_1230, n_6_1229, n_6_1228, n_6_1227, n_6_1226, 
    n_6_1225, n_6_1224, n_6_1223, n_6_1222, n_6_1221, n_6_1220, n_6_1219, n_6_1218, 
    n_6_1217, n_6_1216, n_6_1215}), .Multiplier ({Multiplier[31], hfn_ipo_n27, drc_ipo_n26625, 
    drc_ipo_n26624, drc_ipoPP_7, Multiplier[26], drc_ipo_n26621, drc_ipo_n26620, 
    drc_ipo_n26618, drc_ipo_n26617, drc_ipo_n26616, drc_ipo_n26615, drc_ipo_n26614, 
    drc_ipo_n26613, drc_ipoPP_4, CLOCK_sgo__n46808, drc_ipo_n26610, drc_ipo_n26609, 
    CLOCK_sgo__n46814, drc_ipo_n26607, drc_ipo_n26606, drc_ipo_n26605, drc_ipoPP_1, 
    drc_ipoPP_0, drc_ipo_n26602, drc_ipo_n26599, drc_ipo_n26600, slo__n4944, slo__n3804, 
    sgo__n1306, drc_ipo_n26598, hfn_ipo_n29}), .p_0 ({uc_37, n_6_2354, opt_ipo_n45138, 
    n_6_2352, slo__n18084, n_6_2350, n_6_2349, n_6_2348, CLOCK_slo__n57899, n_6_2346, 
    n_6_2345, n_6_2344, slo__n38018, n_6_2342, n_6_2341, n_6_2340, n_6_2339, slo__n36610, 
    n_6_2337, n_6_2336, n_6_2335, n_6_2334, slo__n17338, slo___n17155, opt_ipo_n23778, 
    slo__n18178, n_6_2329, opt_ipo_n26244, opt_ipo_n24251, slo___n16361, CLOCK_opt_ipo_n45918, 
    n_6_2324}));
datapath__0_187 i_6_75 (.p_2 ({n_6_1214, n_6_1213, n_6_1212, n_6_1211, n_6_1210, 
    n_6_1209, n_6_1208, n_6_1207, n_6_1206, n_6_1205, n_6_1204, n_6_1203, n_6_1202, 
    n_6_1201, n_6_1200, n_6_1199, n_6_1198, n_6_1197, n_6_1196, n_6_1195, n_6_1194, 
    n_6_1193, n_6_1192, n_6_1191, n_6_1190, n_6_1189, n_6_1188, n_6_1187, n_6_1186, 
    n_6_1185, n_6_1184, n_6_1183}), .p_0 ({n_6_30, hfn_ipo_n32, drc_ipo_n26573, drc_ipo_n26574, 
    n_6_26, n_6_25, drc_ipo_n26575, CLOCK_sgo__n47049, drc_ipo_n26576, drc_ipo_n26577, 
    drc_ipo_n26579, drc_ipo_n26581, drc_ipo_n26582, drc_ipo_n26583, drc_ipo_n26585, 
    drc_ipo_n26584, drc_ipo_n26586, drc_ipo_n26587, drc_ipo_n26588, drc_ipo_n26589, 
    drc_ipo_n26592, drc_ipo_n26590, slo__n26645, slo__n4932, slo__n26805, slo__n26713, 
    slo__n16572, slo__n26761, slo__n3800, slo__n16608, slo__n31700, hfn_ipo_n29})
    , .p_1 ({uc_36, opt_ipo_n45145, n_6_2384, n_6_2383, n_6_2382, n_6_2381, n_6_2380, 
    n_6_2379, n_6_2378, n_6_2377, n_6_2376, n_6_2375, n_6_2374, n_6_2373, n_6_2372, 
    n_6_2371, n_6_2370, slo___n19058, slo__n16152, n_6_2367, n_6_2366, slo__n19179, 
    n_6_2364, slo__n30671, n_6_2362, n_6_2361, n_6_2360, n_6_2359, slo___n17582, 
    n_6_2357, n_6_2356, n_6_2355}), .opt_ipoPP_1 (opt_ipo_n45144));
datapath__0_186 i_6_74 (.p_1 ({n_6_1182, n_6_1181, n_6_1180, n_6_1179, n_6_1178, 
    n_6_1177, n_6_1176, n_6_1175, n_6_1174, n_6_1173, n_6_1172, n_6_1171, n_6_1170, 
    n_6_1169, n_6_1168, n_6_1167, n_6_1166, n_6_1165, n_6_1164, n_6_1163, n_6_1162, 
    n_6_1161, n_6_1160, n_6_1159, n_6_1158, n_6_1157, n_6_1156, n_6_1155, n_6_1154, 
    n_6_1153, n_6_1152, n_6_1151}), .Multiplier ({Multiplier[31], hfn_ipo_n27, drc_ipo_n26625, 
    drc_ipo_n26624, drc_ipoPP_7, Multiplier[26], drc_ipo_n26621, drc_ipo_n26620, 
    drc_ipo_n26618, drc_ipo_n26617, drc_ipo_n26616, drc_ipo_n26615, drc_ipo_n26614, 
    drc_ipo_n26613, drc_ipoPP_4, CLOCK_sgo__n46808, drc_ipo_n26610, drc_ipo_n26609, 
    CLOCK_sgo__n46814, drc_ipo_n26607, drc_ipo_n26606, drc_ipo_n26605, drc_ipoPP_1, 
    drc_ipoPP_0, drc_ipo_n26602, drc_ipo_n26599, drc_ipo_n26600, slo__n4944, slo__n3804, 
    sgo__n1306, drc_ipo_n26598, hfn_ipo_n29}), .p_0 ({uc_35, opt_ipo_n45145, n_6_2384, 
    n_6_2383, slo__n17041, n_6_2381, slo__n16267, n_6_2379, n_6_2378, CLOCK_slo__n57874, 
    n_6_2376, n_6_2375, n_6_2374, CLOCK_slo__n55511, n_6_2372, n_6_2371, n_6_2370, 
    slo___n19058, n_6_2368, slo__n16984, n_6_2366, n_6_2365, n_6_2364, slo__n30670, 
    slo__n17399, n_6_2361, n_6_2360, n_6_2359, slo__n10331, slo__n13570, n_6_2356, 
    n_6_2355}), .p_0_8_PP_0 (slo__sro_n36913), .opt_ipoPP_0 (n_6_2375), .opt_ipoPP_2 (opt_ipo_n45144));
datapath__0_182 i_6_71 (.p_2 ({n_6_1150, n_6_1149, n_6_1148, n_6_1147, n_6_1146, 
    n_6_1145, n_6_1144, n_6_1143, n_6_1142, n_6_1141, n_6_1140, n_6_1139, n_6_1138, 
    n_6_1137, n_6_1136, n_6_1135, n_6_1134, n_6_1133, n_6_1132, n_6_1131, n_6_1130, 
    n_6_1129, n_6_1128, n_6_1127, n_6_1126, n_6_1125, n_6_1124, n_6_1123, n_6_1122, 
    n_6_1121, n_6_1120, n_6_1119}), .p_0 ({n_6_30, hfn_ipo_n32, drc_ipo_n26573, drc_ipo_n26574, 
    n_6_26, n_6_25, drc_ipo_n26575, CLOCK_sgo__n47049, drc_ipo_n26576, drc_ipo_n26577, 
    drc_ipo_n26579, drc_ipo_n26581, drc_ipo_n26582, drc_ipo_n26583, drc_ipo_n26585, 
    drc_ipo_n26584, drc_ipo_n26586, drc_ipo_n26587, drc_ipo_n26588, drc_ipo_n26589, 
    drc_ipo_n26592, drc_ipo_n26590, slo__n26645, slo__n4932, slo__n26805, slo__n26713, 
    slo__n16572, slo__n26761, slo__n3800, slo__n16608, slo__n31700, hfn_ipo_n29})
    , .p_1 ({uc_34, n_6_2416, n_6_2415, n_6_2414, n_6_2413, CLOCK_slo__n55287, n_6_2411, 
    n_6_2410, n_6_2409, n_6_2408, n_6_1_542, n_6_2406, n_6_2405, n_6_2404, n_6_2403, 
    n_6_2402, slo__n16975, slo___n15030, slo__n35114, n_6_2398, n_6_2397, slo__sro_n7405, 
    n_6_2395, slo__n13501, n_6_2393, n_6_2392, n_6_2391, n_6_2390, slo___n6965, CLOCK_opt_ipo_n45825, 
    slo___n7115, n_6_2386}));
datapath__0_181 i_6_70 (.p_1 ({n_6_1118, n_6_1117, n_6_1116, n_6_1115, n_6_1114, 
    n_6_1113, n_6_1112, n_6_1111, n_6_1110, n_6_1109, n_6_1108, n_6_1107, n_6_1106, 
    n_6_1105, n_6_1104, n_6_1103, n_6_1102, n_6_1101, n_6_1100, n_6_1099, n_6_1098, 
    n_6_1097, n_6_1096, n_6_1095, n_6_1094, n_6_1093, n_6_1092, n_6_1091, n_6_1090, 
    n_6_1089, n_6_1088, n_6_1087}), .Multiplier ({Multiplier[31], hfn_ipo_n27, drc_ipo_n26625, 
    drc_ipo_n26624, drc_ipoPP_7, Multiplier[26], drc_ipo_n26621, drc_ipo_n26620, 
    drc_ipo_n26618, drc_ipo_n26617, drc_ipo_n26616, drc_ipo_n26615, drc_ipo_n26614, 
    drc_ipo_n26613, drc_ipoPP_4, CLOCK_sgo__n46808, drc_ipo_n26610, drc_ipo_n26609, 
    CLOCK_sgo__n46814, drc_ipo_n26607, drc_ipo_n26606, drc_ipo_n26605, drc_ipoPP_1, 
    drc_ipoPP_0, drc_ipo_n26602, drc_ipo_n26599, drc_ipo_n26600, slo__n4944, slo__n3804, 
    sgo__n1306, drc_ipo_n26598, hfn_ipo_n29}), .p_0 ({uc_33, n_6_2416, n_6_2415, 
    slo__n17214, n_6_2413, n_6_2412, n_6_2411, n_6_2410, slo__n14465, n_6_2408, n_6_1_542, 
    n_6_2406, CLOCK_slo__n57906, n_6_2404, n_6_2403, n_6_2402, n_6_2401, slo__n11164, 
    slo__n35114, n_6_2398, n_6_2397, slo__sro_n7405, n_6_2395, n_6_2394, n_6_2393, 
    n_6_2392, n_6_2391, n_6_2390, slo___n6965, CLOCK_opt_ipo_n45825, slo___n7115, 
    n_6_2386}));
datapath__0_177 i_6_67 (.p_2 ({n_6_1086, n_6_1085, n_6_1084, n_6_1083, n_6_1082, 
    n_6_1081, n_6_1080, n_6_1079, n_6_1078, n_6_1077, n_6_1076, n_6_1075, n_6_1074, 
    n_6_1073, n_6_1072, n_6_1071, n_6_1070, n_6_1069, n_6_1068, n_6_1067, n_6_1066, 
    n_6_1065, n_6_1064, n_6_1063, n_6_1062, n_6_1061, n_6_1060, n_6_1059, n_6_1058, 
    n_6_1057, n_6_1056, n_6_1055}), .p_0 ({n_6_30, hfn_ipo_n31, drc_ipo_n26573, drc_ipo_n26574, 
    n_6_26, n_6_25, drc_ipo_n26575, CLOCK_sgo__n47049, drc_ipo_n26576, drc_ipo_n26577, 
    drc_ipo_n26579, drc_ipo_n26581, drc_ipo_n26582, drc_ipo_n26583, drc_ipo_n26585, 
    drc_ipo_n26584, drc_ipo_n26586, drc_ipo_n26587, drc_ipo_n26588, drc_ipo_n26589, 
    drc_ipo_n26592, drc_ipo_n26590, slo__n26645, slo__n4932, slo__n26805, slo__n26713, 
    slo__n16572, slo__n26761, slo__n3800, slo__n16608, slo__n31700, hfn_ipo_n29})
    , .p_1 ({uc_32, n_6_2447, n_6_2446, opt_ipo_n24966, n_6_2444, slo__sro_n8179, 
    n_6_2442, opt_ipo_n24743, n_6_2440, n_6_2439, n_6_2438, n_6_2437, n_6_2436, n_6_2435, 
    opt_ipo_n24861, n_6_2433, n_6_2432, n_6_2431, n_6_2430, n_6_2429, CLOCK_opt_ipo_n46005, 
    slo__n35802, n_6_2426, slo__n11420, n_6_2424, n_6_2423, slo__n18523, n_6_2421, 
    n_6_2420, n_6_2419, n_6_2418, n_6_2417}));
datapath__0_176 i_6_66 (.p_1 ({n_6_1054, n_6_1053, n_6_1052, n_6_1051, n_6_1050, 
    n_6_1049, n_6_1048, n_6_1047, n_6_1046, n_6_1045, n_6_1044, n_6_1043, n_6_1042, 
    n_6_1041, n_6_1040, n_6_1039, n_6_1038, n_6_1037, n_6_1036, n_6_1035, n_6_1034, 
    n_6_1033, n_6_1032, n_6_1031, n_6_1030, n_6_1029, n_6_1028, n_6_1027, n_6_1026, 
    n_6_1025, n_6_1024, n_6_1023}), .Multiplier ({Multiplier[31], hfn_ipo_n26, drc_ipo_n26625, 
    drc_ipo_n26624, drc_ipoPP_7, Multiplier[26], drc_ipo_n26621, drc_ipo_n26620, 
    drc_ipo_n26618, drc_ipo_n26617, drc_ipo_n26616, drc_ipo_n26615, drc_ipo_n26614, 
    drc_ipo_n26613, drc_ipoPP_4, CLOCK_sgo__n46808, drc_ipo_n26610, drc_ipo_n26609, 
    CLOCK_sgo__n46814, drc_ipo_n26607, drc_ipo_n26606, drc_ipo_n26605, drc_ipoPP_1, 
    drc_ipoPP_0, drc_ipo_n26602, drc_ipo_n26599, drc_ipo_n26600, slo__n4944, slo__n3804, 
    sgo__n1306, drc_ipo_n26598, hfn_ipo_n29}), .p_0 ({uc_31, n_6_2447, n_6_2446, 
    opt_ipo_n24966, n_6_2444, slo__sro_n8179, n_6_2442, opt_ipo_n24743, CLOCK_slo__n53562, 
    n_6_2439, n_6_2438, n_6_2437, slo__n17575, n_6_2435, opt_ipo_n24861, n_6_2433, 
    n_6_2432, n_6_2431, n_6_2430, slo__n12976, CLOCK_opt_ipo_n46005, slo__n35802, 
    n_6_2426, n_6_2425, slo__n18286, n_6_2423, n_6_2422, n_6_2421, n_6_2420, n_6_2419, 
    n_6_2418, n_6_2417}));
datapath__0_172 i_6_63 (.p_2 ({n_6_1022, n_6_1021, n_6_1020, n_6_1019, n_6_1018, 
    n_6_1017, n_6_1016, n_6_1015, n_6_1014, n_6_1013, n_6_1012, n_6_1011, n_6_1010, 
    n_6_1009, n_6_1008, n_6_1007, n_6_1006, n_6_1005, n_6_1004, n_6_1003, n_6_1002, 
    n_6_1001, n_6_1000, n_6_999, n_6_998, n_6_997, n_6_996, n_6_995, n_6_994, n_6_993, 
    n_6_992, n_6_991}), .p_0 ({n_6_30, hfn_ipo_n31, drc_ipo_n26573, drc_ipo_n26574, 
    n_6_26, n_6_25, drc_ipo_n26575, CLOCK_sgo__n47049, drc_ipo_n26576, drc_ipo_n26577, 
    drc_ipo_n26579, drc_ipo_n26581, drc_ipo_n26582, drc_ipo_n26583, drc_ipo_n26585, 
    drc_ipo_n26584, drc_ipo_n26586, drc_ipo_n26587, drc_ipo_n26588, drc_ipo_n26589, 
    drc_ipo_n26592, drc_ipo_n26590, slo__n26645, slo__n4932, slo__n26805, slo__n26713, 
    slo__n16572, slo__n26761, slo__n3800, slo__n16608, slo__n31700, hfn_ipo_n29})
    , .p_1 ({uc_30, n_6_2478, n_6_2477, n_6_2476, n_6_2475, n_6_2474, opt_ipo_n45366, 
    n_6_2472, n_6_2471, n_6_2470, n_6_2469, n_6_2468, n_6_2467, n_6_2466, n_6_2465, 
    n_6_2464, n_6_2463, n_6_2462, n_6_2461, n_6_2460, n_6_2459, opt_ipo_n25394, n_6_2457, 
    n_6_2456, n_6_2455, slo___n17886, slo__n13417, n_6_2452, n_6_2451, n_6_2450, 
    slo__n31336, n_6_2448}));
datapath__0_171 i_6_62 (.p_1 ({n_6_990, n_6_989, n_6_988, n_6_987, n_6_986, n_6_985, 
    n_6_984, n_6_983, n_6_982, n_6_981, n_6_980, n_6_979, n_6_978, n_6_977, n_6_976, 
    n_6_975, n_6_974, n_6_973, n_6_972, n_6_971, n_6_970, n_6_969, n_6_968, n_6_967, 
    n_6_966, n_6_965, n_6_964, n_6_963, n_6_962, n_6_961, n_6_960, n_6_959}), .Multiplier ({
    Multiplier[31], hfn_ipo_n26, drc_ipo_n26625, drc_ipo_n26624, drc_ipoPP_7, Multiplier[26], 
    drc_ipo_n26621, drc_ipo_n26620, drc_ipo_n26618, drc_ipo_n26617, drc_ipo_n26616, 
    drc_ipo_n26615, drc_ipo_n26614, drc_ipo_n26613, drc_ipoPP_4, CLOCK_sgo__n46808, 
    drc_ipo_n26610, drc_ipo_n26609, CLOCK_sgo__n46814, drc_ipo_n26607, drc_ipo_n26606, 
    drc_ipo_n26605, drc_ipoPP_1, drc_ipoPP_0, drc_ipo_n26602, drc_ipo_n26599, drc_ipo_n26600, 
    slo__n4944, slo__n3804, sgo__n1306, drc_ipo_n26598, hfn_ipo_n29}), .p_0 ({uc_29, 
    n_6_2478, n_6_2477, n_6_2476, n_6_2475, n_6_2474, opt_ipo_n45366, CLOCK_slo__n54964, 
    n_6_2471, n_6_2470, n_6_2469, n_6_2468, n_6_2467, n_6_2466, n_6_2465, slo__n14037, 
    slo__n16706, n_6_2462, n_6_2461, n_6_2460, n_6_2459, opt_ipo_n25394, n_6_2457, 
    n_6_2456, n_6_2455, slo___n17886, n_6_2453, n_6_2452, slo__n17744, n_6_2450, 
    slo__n31336, n_6_2448}));
datapath__0_167 i_6_59 (.p_2 ({n_6_958, n_6_957, n_6_956, n_6_955, n_6_954, n_6_953, 
    n_6_952, n_6_951, n_6_950, n_6_949, n_6_948, n_6_947, n_6_946, n_6_945, n_6_944, 
    n_6_943, n_6_942, n_6_941, n_6_940, n_6_939, n_6_938, n_6_937, n_6_936, n_6_935, 
    n_6_934, n_6_933, n_6_932, n_6_931, n_6_930, n_6_929, n_6_928, n_6_927}), .p_0 ({
    n_6_30, hfn_ipo_n31, drc_ipo_n26573, drc_ipo_n26574, n_6_26, n_6_25, drc_ipo_n26575, 
    CLOCK_sgo__n47049, drc_ipo_n26576, drc_ipo_n26577, drc_ipo_n26579, n_6_19, drc_ipo_n26582, 
    drc_ipo_n26583, drc_ipo_n26585, drc_ipo_n26584, drc_ipo_n26586, drc_ipo_n26587, 
    drc_ipo_n26588, drc_ipo_n26589, drc_ipo_n26592, drc_ipo_n26590, slo__n26645, 
    slo__n4932, slo__n26805, slo__n26713, slo__n16572, slo__n26761, slo__n3800, slo__n16608, 
    slo__n31700, hfn_ipo_n29}), .p_1 ({uc_28, n_6_2509, n_6_2508, n_6_2507, n_6_2506, 
    n_6_2505, n_6_2504, n_6_2503, n_6_2502, n_6_2501, n_6_2500, slo__n13621, n_6_2498, 
    n_6_2497, n_6_2496, n_6_2495, n_6_2494, n_6_2493, n_6_2492, n_6_2491, n_6_2490, 
    n_6_2489, n_6_2488, n_6_2487, n_6_2486, slo__n14026, slo__n13938, slo__n14126, 
    n_6_2482, slo__n13933, slo__n14113, n_6_2479}));
datapath__0_166 i_6_58 (.p_1 ({n_6_926, n_6_925, n_6_924, n_6_923, n_6_922, n_6_921, 
    n_6_920, n_6_919, n_6_918, n_6_917, n_6_916, n_6_915, n_6_914, n_6_913, n_6_912, 
    n_6_911, n_6_910, n_6_909, n_6_908, n_6_907, n_6_906, n_6_905, n_6_904, n_6_903, 
    n_6_902, n_6_901, n_6_900, n_6_899, n_6_898, n_6_897, n_6_896, n_6_895}), .Multiplier ({
    Multiplier[31], hfn_ipo_n26, drc_ipo_n26625, drc_ipo_n26624, drc_ipoPP_7, Multiplier[26], 
    drc_ipo_n26621, drc_ipo_n26620, drc_ipo_n26618, drc_ipo_n26617, drc_ipo_n26616, 
    drc_ipo_n26615, drc_ipo_n26614, drc_ipo_n26613, drc_ipoPP_4, CLOCK_sgo__n46808, 
    drc_ipo_n26610, drc_ipo_n26609, CLOCK_sgo__n46814, drc_ipo_n26607, Multiplier[11], 
    drc_ipo_n26605, drc_ipoPP_1, drc_ipoPP_0, drc_ipo_n26602, drc_ipo_n26599, drc_ipo_n26600, 
    slo__n4944, slo__n3804, sgo__n1306, drc_ipo_n26598, hfn_ipo_n29}), .p_0 ({uc_27, 
    n_6_2509, n_6_2508, n_6_2507, n_6_2506, n_6_2505, slo__n12811, n_6_2503, slo__n12606, 
    n_6_2501, n_6_2500, n_6_2499, n_6_2498, n_6_2497, n_6_2496, n_6_2495, n_6_2494, 
    slo__n38401, n_6_2492, n_6_2491, n_6_2490, CLOCK_slo__n53697, n_6_2488, n_6_2487, 
    n_6_2486, n_6_2485, n_6_2484, n_6_2483, n_6_2482, n_6_2481, n_6_2480, n_6_2479})
    , .drc_ipoPP_0 (drc_ipo_n26606));
datapath__0_162 i_6_55 (.p_2 ({n_6_894, n_6_893, n_6_892, n_6_891, n_6_890, n_6_889, 
    n_6_888, n_6_887, n_6_886, n_6_885, n_6_884, n_6_883, n_6_882, n_6_881, n_6_880, 
    n_6_879, n_6_878, n_6_877, n_6_876, n_6_875, n_6_874, n_6_873, n_6_872, n_6_871, 
    n_6_870, n_6_869, n_6_868, n_6_867, n_6_866, n_6_865, n_6_864, n_6_863}), .p_0 ({
    n_6_30, hfn_ipo_n31, drc_ipo_n26573, drc_ipo_n26574, n_6_26, n_6_25, drc_ipo_n26575, 
    CLOCK_sgo__n47049, drc_ipo_n26576, n_6_21, drc_ipo_n26579, n_6_19, CLOCK_sgo__n47026, 
    drc_ipo_n26583, n_6_16, n_6_15, drc_ipo_n26586, drc_ipo_n26587, n_6_12, drc_ipo_n26589, 
    drc_ipo_n26592, drc_ipo_n26591, slo__n26645, slo__n4932, slo__n26805, slo__n26713, 
    slo__n16572, slo__n26761, slo__n3800, slo__n16608, slo__n31700, hfn_ipo_n29})
    , .p_1 ({uc_26, n_6_2540, n_6_2539, n_6_2538, n_6_2537, slo___n9717, n_6_2535, 
    n_6_2534, slo__n13610, n_6_2532, n_6_2531, n_6_2530, n_6_2529, n_6_2528, n_6_2527, 
    n_6_2526, slo__n17556, n_6_2524, n_6_2523, slo___n17357, opt_ipo_n23804, n_6_2520, 
    n_6_2519, n_6_2518, n_6_2517, slo___n6972, CLOCK_slo___n52225, n_6_2514, n_6_2513, 
    opt_ipo_n24285, n_6_2511, n_6_2510}), .drc_ipoPP_0 (drc_ipo_n26577), .p_0_19_PP_0 (CLOCK_sgo__n47026));
datapath__0_161 i_6_54 (.p_1 ({n_6_862, n_6_861, n_6_860, n_6_859, n_6_858, n_6_857, 
    n_6_856, n_6_855, n_6_854, n_6_853, n_6_852, n_6_851, n_6_850, n_6_849, n_6_848, 
    n_6_847, n_6_846, n_6_845, n_6_844, n_6_843, n_6_842, n_6_841, n_6_840, n_6_839, 
    n_6_838, n_6_837, n_6_836, n_6_835, n_6_834, n_6_833, n_6_832, n_6_831}), .Multiplier ({
    Multiplier[31], hfn_ipo_n26, drc_ipo_n26625, drc_ipo_n26624, drc_ipoPP_7, Multiplier[26], 
    drc_ipo_n26621, drc_ipo_n26620, drc_ipoPP_5, drc_ipo_n26617, drc_ipo_n26616, 
    drc_ipo_n26615, CLOCK_sgo__n46725, drc_ipo_n26613, drc_ipoPP_4, CLOCK_sgo__n46808, 
    drc_ipo_n26610, drc_ipo_n26609, CLOCK_sgo__n46815, drc_ipo_n26607, Multiplier[11], 
    drc_ipo_n26605, drc_ipoPP_1, drc_ipoPP_0, drc_ipo_n26602, drc_ipo_n26599, drc_ipo_n26600, 
    slo__n4944, slo__n3804, sgo__n1306, drc_ipo_n26598, hfn_ipo_n29}), .p_0 ({uc_25, 
    n_6_2540, n_6_2539, n_6_2538, n_6_2537, slo___n9717, n_6_2535, n_6_2534, n_6_2533, 
    CLOCK_slo__n56953, CLOCK_slo__n56933, n_6_2530, n_6_2529, n_6_2528, slo__n16871, 
    slo__n39136, n_6_2525, n_6_2524, n_6_2523, slo__n11427, opt_ipo_n23804, n_6_2520, 
    n_6_2519, n_6_2518, n_6_2517, slo___n6972, CLOCK_slo___n52225, n_6_2514, n_6_2513, 
    opt_ipo_n24285, n_6_2511, n_6_2510}), .drc_ipoPP_0 (drc_ipo_n26614));
datapath__0_157 i_6_51 (.p_2 ({n_6_830, n_6_829, n_6_828, n_6_827, n_6_826, n_6_825, 
    n_6_824, n_6_823, n_6_822, n_6_821, n_6_820, n_6_819, n_6_818, n_6_817, n_6_816, 
    n_6_815, n_6_814, n_6_813, n_6_812, n_6_811, n_6_810, n_6_809, n_6_808, n_6_807, 
    n_6_806, n_6_805, n_6_804, n_6_803, n_6_802, n_6_801, n_6_800, n_6_799}), .p_0 ({
    n_6_30, hfn_ipo_n31, n_6_28, drc_ipo_n26574, n_6_26, n_6_25, drc_ipo_n26575, 
    CLOCK_sgo__n47050, n_6_22, n_6_21, n_6_20, n_6_19, CLOCK_sgo__n47026, n_6_17, 
    n_6_16, n_6_15, drc_ipo_n26586, drc_ipo_n26587, n_6_12, n_6_11, n_6_10, drc_ipo_n26591, 
    slo__n26645, slo__n4932, slo__n26805, slo__n26713, slo__n16572, slo__n26761, 
    slo__n3800, slo__n16608, slo__n31700, hfn_ipo_n29}), .p_1 ({uc_24, n_6_2571, 
    n_6_2570, n_6_2569, n_6_2568, n_6_2567, n_6_2566, n_6_2565, n_6_2564, n_6_2563, 
    n_6_2562, n_6_2561, n_6_2560, n_6_2559, n_6_2558, n_6_2557, slo__n14709, n_6_2555, 
    n_6_2554, slo__n14696, n_6_2552, n_6_2551, slo__n14899, n_6_2549, n_6_2548, n_6_2547, 
    n_6_2546, n_6_2545, slo__n14062, slo__n14691, n_6_2542, n_6_2541}));
datapath__0_156 i_6_50 (.p_1 ({n_6_798, n_6_797, n_6_796, n_6_795, n_6_794, n_6_793, 
    n_6_792, n_6_791, n_6_790, n_6_789, n_6_788, n_6_787, n_6_786, n_6_785, n_6_784, 
    n_6_783, n_6_782, n_6_781, n_6_780, n_6_779, n_6_778, n_6_777, n_6_776, n_6_775, 
    n_6_774, n_6_773, n_6_772, n_6_771, n_6_770, n_6_769, n_6_768, n_6_767}), .Multiplier ({
    Multiplier[31], hfn_ipo_n26, drc_ipo_n26625, drc_ipo_n26624, drc_ipoPP_7, drc_ipoPP_6, 
    drc_ipo_n26621, drc_ipo_n26620, drc_ipoPP_5, drc_ipo_n26617, Multiplier[21], 
    drc_ipo_n26615, CLOCK_sgo__n46725, drc_ipo_n26613, drc_ipoPP_4, CLOCK_sgo__n46808, 
    Multiplier[15], drc_ipo_n26609, CLOCK_sgo__n46815, Multiplier[12], Multiplier[11], 
    drc_ipo_n26605, drc_ipoPP_1, drc_ipoPP_0, drc_ipo_n26602, drc_ipo_n26599, drc_ipo_n26600, 
    slo__n4944, slo__n3804, sgo__n1306, drc_ipo_n26598, hfn_ipo_n29}), .p_0 ({uc_23, 
    n_6_2571, n_6_2570, n_6_2569, n_6_2568, CLOCK_slo__n56237, n_6_2566, n_6_2565, 
    CLOCK_slo__n56946, n_6_2563, slo__n16343, n_6_2561, n_6_2560, n_6_2559, n_6_2558, 
    slo__n19255, n_6_2556, n_6_2555, n_6_2554, n_6_2553, n_6_2552, slo__n18942, slo___n17474, 
    n_6_2549, slo__n18973, n_6_2547, n_6_2546, n_6_2545, n_6_2544, n_6_2543, slo__n12071, 
    n_6_2541}));
datapath__0_152 i_6_47 (.p_2 ({n_6_766, n_6_765, n_6_764, n_6_763, n_6_762, n_6_761, 
    n_6_760, n_6_759, n_6_758, n_6_757, n_6_756, n_6_755, n_6_754, n_6_753, n_6_752, 
    n_6_751, n_6_750, n_6_749, n_6_748, n_6_747, n_6_746, n_6_745, n_6_744, n_6_743, 
    n_6_742, n_6_741, n_6_740, n_6_739, n_6_738, n_6_737, n_6_736, n_6_735}), .p_0 ({
    n_6_30, hfn_ipo_n31, n_6_28, drc_ipo_n26574, n_6_26, n_6_25, drc_ipo_n26575, 
    CLOCK_sgo__n47050, n_6_22, n_6_21, n_6_20, n_6_19, CLOCK_sgo__n47026, n_6_17, 
    n_6_16, n_6_15, n_6_14, n_6_13, n_6_12, n_6_11, n_6_10, drc_ipo_n26591, slo__n26648, 
    slo__n4932, slo__n26805, slo__n26713, slo__n16572, slo__n26761, slo__n3800, slo__n16608, 
    slo__n31700, hfn_ipo_n29}), .p_1 ({uc_22, n_6_2602, n_6_2601, n_6_2600, slo__n35732, 
    n_6_1_757, n_6_2597, n_6_2596, n_6_2595, n_6_2594, n_6_2593, n_6_2592, n_6_2591, 
    n_6_2590, n_6_2589, n_6_2588, slo__n14942, n_6_2586, n_6_2585, n_6_2584, n_6_2583, 
    n_6_2582, n_6_2581, CLOCK_opt_ipo_n46029, slo__n12190, opt_ipo_n44599, slo__n37437, 
    n_6_2576, n_6_1_734, n_6_2574, n_6_2573, spw__n67889}));
datapath__0_151 i_6_46 (.p_1 ({n_6_734, n_6_733, n_6_732, n_6_731, n_6_730, n_6_729, 
    n_6_728, n_6_727, n_6_726, n_6_725, n_6_724, n_6_723, n_6_722, n_6_721, n_6_720, 
    n_6_719, n_6_718, n_6_717, n_6_716, n_6_715, n_6_714, n_6_713, n_6_712, n_6_711, 
    n_6_710, n_6_709, n_6_708, n_6_707, n_6_706, n_6_705, n_6_704, n_6_703}), .Multiplier ({
    Multiplier[31], hfn_ipo_n26, Multiplier[29], drc_ipo_n26624, drc_ipoPP_7, drc_ipoPP_6, 
    CLOCK_sgo__n46841, drc_ipo_n26620, drc_ipoPP_5, drc_ipo_n26617, Multiplier[21], 
    drc_ipo_n26615, CLOCK_sgo__n46725, Multiplier[18], drc_ipoPP_4, drc_ipoPP_3PP_0, 
    Multiplier[15], drc_ipo_n26609, CLOCK_sgo__n46815, Multiplier[12], Multiplier[11], 
    drc_ipo_n26605, drc_ipoPP_1, drc_ipoPP_0, drc_ipo_n26602, drc_ipo_n26599, drc_ipo_n26600, 
    slo__n4944, slo__n3804, sgo__n1306, drc_ipo_n26598, hfn_ipo_n29}), .p_0 ({uc_21, 
    n_6_2602, slo__n10168, n_6_2600, slo__n35732, n_6_1_757, slo__n14486, n_6_2596, 
    n_6_2595, n_6_2594, CLOCK_slo__n56232, n_6_2592, n_6_2591, n_6_2590, n_6_2589, 
    n_6_2588, n_6_2587, n_6_2586, n_6_2585, n_6_2584, n_6_2583, n_6_2582, slo__n37202, 
    CLOCK_opt_ipo_n46029, slo___n13777, opt_ipo_n44599, n_6_2577, n_6_2576, n_6_1_734, 
    n_6_2574, n_6_2573, spw__n67889}));
datapath__0_147 i_6_43 (.p_2 ({n_6_702, n_6_701, n_6_700, n_6_699, n_6_698, n_6_697, 
    n_6_696, n_6_695, n_6_694, n_6_693, n_6_692, n_6_691, n_6_690, n_6_689, n_6_688, 
    n_6_687, n_6_686, n_6_685, n_6_684, n_6_683, n_6_682, n_6_681, n_6_680, n_6_679, 
    n_6_678, n_6_677, n_6_676, n_6_675, n_6_674, n_6_673, n_6_672, n_6_671}), .p_0 ({
    n_6_30, hfn_ipo_n31, n_6_28, drc_ipo_n26574, n_6_26, n_6_25, drc_ipo_n26575, 
    CLOCK_sgo__n47050, n_6_22, n_6_21, n_6_20, n_6_19, CLOCK_sgo__n47026, n_6_17, 
    n_6_16, n_6_15, n_6_14, n_6_13, n_6_12, n_6_11, n_6_10, drc_ipo_n26591, slo__n26648, 
    slo__n4932, slo__n26805, slo__n26713, slo__n16572, slo__n26761, slo__n3800, slo__n16608, 
    slo__n31700, sgo__n1276}), .p_1 ({uc_20, n_6_2633, n_6_2632, n_6_2631, n_6_2630, 
    n_6_2629, n_6_2628, n_6_2627, n_6_2626, n_6_2625, slo___n12846, n_6_2623, n_6_2622, 
    n_6_2621, opt_ipo_n24166, n_6_1_782, n_6_2618, n_6_2617, slo__n37463, slo__n38656, 
    n_6_2614, n_6_2613, n_6_2612, n_6_2611, n_6_2610, n_6_2609, n_6_2608, n_6_2607, 
    CLOCK_slo__sro_n58313, CLOCK_slo___n54911, n_6_2604, CLOCK_slo___n64354}), .opt_ipoPP_1 (opt_ipo_n44394));
datapath__0_146 i_6_42 (.p_1 ({n_6_670, n_6_669, n_6_668, n_6_667, n_6_666, n_6_665, 
    n_6_664, n_6_663, n_6_662, n_6_661, n_6_660, n_6_659, n_6_658, n_6_657, n_6_656, 
    n_6_655, n_6_654, n_6_653, n_6_652, n_6_651, n_6_650, n_6_649, n_6_648, n_6_647, 
    n_6_646, n_6_645, n_6_644, n_6_643, n_6_642, n_6_641, n_6_640, n_6_639}), .Multiplier ({
    Multiplier[31], hfn_ipo_n26, Multiplier[29], drc_ipo_n26624, Multiplier[27], 
    drc_ipoPP_6, CLOCK_sgo__n46841, drc_ipo_n26620, drc_ipoPP_5, drc_ipo_n26617, 
    Multiplier[21], drc_ipo_n26615, CLOCK_sgo__n46725, Multiplier[18], drc_ipoPP_4, 
    drc_ipoPP_3, Multiplier[15], drc_ipo_n26609, CLOCK_sgo__n46815, Multiplier[12], 
    Multiplier[11], drc_ipo_n26605, drc_ipoPP_1, drc_ipoPP_0, drc_ipo_n26602, drc_ipo_n26599, 
    drc_ipo_n26600, slo__n4944, slo__n3804, sgo__n1306, drc_ipo_n26598, sgo__n1276})
    , .p_0 ({uc_19, n_6_2633, n_6_2632, n_6_2631, n_6_2630, CLOCK_slo__n55647, slo__n7753, 
    n_6_2627, slo__n11270, n_6_2625, slo___n12846, n_6_2623, CLOCK_slo__n57518, n_6_2621, 
    CLOCK_slo__n57547, n_6_1_782, n_6_2618, n_6_2617, n_6_2616, n_6_2615, slo__n13910, 
    slo__n37415, n_6_2612, n_6_2611, n_6_2610, slo__n38227, n_6_2608, n_6_2607, CLOCK_slo__sro_n58313, 
    CLOCK_slo___n54911, n_6_2604, CLOCK_slo___n64354}), .opt_ipoPP_1 (opt_ipo_n44394));
datapath__0_142 i_6_39 (.p_2 ({n_6_638, n_6_637, n_6_636, n_6_635, n_6_634, n_6_633, 
    n_6_632, n_6_631, n_6_630, n_6_629, n_6_628, n_6_627, n_6_626, n_6_625, n_6_624, 
    n_6_623, n_6_622, n_6_621, n_6_620, n_6_619, n_6_618, n_6_617, n_6_616, n_6_615, 
    n_6_614, n_6_613, n_6_612, n_6_611, n_6_610, n_6_609, n_6_608, n_6_607}), .p_0 ({
    n_6_30, hfn_ipo_n30, n_6_28, drc_ipo_n26574, n_6_26, n_6_25, CLOCK_sgo__n47054, 
    CLOCK_sgo__n47050, n_6_22, n_6_21, n_6_20, n_6_19, CLOCK_sgo__n47026, n_6_17, 
    n_6_16, n_6_15, n_6_14, n_6_13, n_6_12, n_6_11, n_6_10, drc_ipo_n26591, slo__n26648, 
    slo__n4932, slo__n26805, slo__n26713, slo__n16572, slo__n26761, slo__n3800, slo__n16608, 
    slo__n31700, sgo__n1276}), .p_1 ({uc_18, n_6_2664, n_6_2663, n_6_2662, n_6_2661, 
    slo__n16796, n_6_2659, CLOCK_slo__n55232, n_6_2657, n_6_2656, slo___n19273, slo___n19182, 
    n_6_2653, slo__n19102, n_6_2651, slo__n19282, n_6_2649, n_6_2648, n_6_2647, n_6_2646, 
    CLOCK_slo__n57556, slo__n13438, slo__n13903, n_6_2642, n_6_2641, n_6_2640, n_6_2639, 
    slo__n36492, slo__n38056, n_6_2636, slo__n11048, n_6_2634}));
datapath__0_141 i_6_38 (.p_1 ({n_6_606, n_6_605, n_6_604, n_6_603, n_6_602, n_6_601, 
    n_6_600, n_6_599, n_6_598, n_6_597, n_6_596, n_6_595, n_6_594, n_6_593, n_6_592, 
    n_6_591, n_6_590, n_6_589, n_6_588, n_6_587, n_6_586, n_6_585, n_6_584, n_6_583, 
    n_6_582, n_6_581, n_6_580, n_6_579, n_6_578, n_6_577, n_6_576, n_6_575}), .Multiplier ({
    Multiplier[31], hfn_ipo_n25, Multiplier[29], drc_ipo_n26624, Multiplier[27], 
    drc_ipoPP_6, CLOCK_sgo__n46841, drc_ipo_n26620, drc_ipoPP_5, drc_ipo_n26617, 
    Multiplier[21], drc_ipo_n26615, CLOCK_sgo__n46725, Multiplier[18], drc_ipoPP_4, 
    drc_ipoPP_3, Multiplier[15], drc_ipo_n26609, CLOCK_sgo__n46815, Multiplier[12], 
    Multiplier[11], drc_ipo_n26605, drc_ipoPP_1, drc_ipoPP_0, drc_ipo_n26602, drc_ipo_n26599, 
    drc_ipo_n26600, slo__n4944, slo__n3804, sgo__n1306, drc_ipo_n26598, sgo__n1276})
    , .p_0 ({uc_17, n_6_2664, n_6_2663, n_6_2662, slo__n16392, n_6_2660, slo__n16413, 
    slo__n16280, slo__n12818, n_6_2656, slo___n19273, slo___n19182, n_6_2653, n_6_2652, 
    n_6_2651, n_6_2650, n_6_2649, n_6_2648, n_6_2647, n_6_2646, n_6_2645, n_6_2644, 
    slo___n15116, n_6_2642, n_6_2641, n_6_2640, n_6_2639, n_6_2638, n_6_2637, n_6_2636, 
    n_6_2635, n_6_2634}));
datapath__0_137 i_6_35 (.p_2 ({n_6_574, n_6_573, n_6_572, n_6_571, n_6_570, n_6_569, 
    n_6_568, n_6_567, n_6_566, n_6_565, n_6_564, n_6_563, n_6_562, n_6_561, n_6_560, 
    n_6_559, n_6_558, n_6_557, n_6_556, n_6_555, n_6_554, n_6_553, n_6_552, n_6_551, 
    n_6_550, n_6_549, n_6_548, n_6_547, n_6_546, n_6_545, n_6_544, n_6_543}), .p_0 ({
    n_6_30, hfn_ipo_n30, n_6_28, drc_ipo_n26574, n_6_26, n_6_25, CLOCK_sgo__n47054, 
    CLOCK_sgo__n47050, n_6_22, n_6_21, n_6_20, n_6_19, CLOCK_sgo__n47026, n_6_17, 
    n_6_16, n_6_15, n_6_14, n_6_13, n_6_12, n_6_11, n_6_10, drc_ipo_n26591, slo__n26654, 
    slo__n4932, slo__n26805, slo__n26713, slo__n16572, slo__n26761, slo__n3800, slo__n16608, 
    slo__n31700, sgo__n1276}), .p_1 ({uc_16, n_6_2695, n_6_2694, slo__n14949, n_6_2692, 
    opt_ipo_n44105, n_6_2690, n_6_2689, n_6_2688, slo__n26895, n_6_2686, n_6_2685, 
    n_6_2684, n_6_2683, n_6_2682, n_6_2681, n_6_2680, slo__n13838, n_6_2678, n_6_2677, 
    n_6_2676, n_6_2675, CLOCK_opt_ipo_n46038, n_6_2673, n_6_2672, slo__sro_n6239, 
    n_6_2670, slo__sro_n15108, n_6_2668, n_6_2667, n_6_2666, n_6_2665}), .p_0_9_PP_0 (slo__n26654));
datapath__0_136 i_6_34 (.p_1 ({n_6_542, n_6_541, n_6_540, n_6_539, n_6_538, n_6_537, 
    n_6_536, n_6_535, n_6_534, n_6_533, n_6_532, n_6_531, n_6_530, n_6_529, n_6_528, 
    n_6_527, n_6_526, n_6_525, n_6_524, n_6_523, n_6_522, n_6_521, n_6_520, n_6_519, 
    n_6_518, n_6_517, n_6_516, n_6_515, n_6_514, n_6_513, n_6_512, n_6_511}), .Multiplier ({
    Multiplier[31], hfn_ipo_n25, Multiplier[29], drc_ipo_n26624, Multiplier[27], 
    drc_ipoPP_6, CLOCK_sgo__n46841, drc_ipo_n26620, drc_ipoPP_5, drc_ipo_n26617, 
    Multiplier[21], drc_ipo_n26615, CLOCK_sgo__n46725, Multiplier[18], drc_ipoPP_4, 
    drc_ipoPP_3, Multiplier[15], drc_ipo_n26609, CLOCK_sgo__n46815, Multiplier[12], 
    Multiplier[11], drc_ipo_n26605, drc_ipoPP_1, drc_ipoPP_0, drc_ipo_n26602, drc_ipo_n26599, 
    drc_ipo_n26600, slo__n4944, slo__n3804, sgo__n1306, drc_ipo_n26598, sgo__n1276})
    , .p_0 ({uc_15, n_6_2695, n_6_2694, n_6_2693, CLOCK_slo__n55908, opt_ipo_n44105, 
    slo__n12473, n_6_2689, n_6_2688, slo__n26894, n_6_2686, n_6_2685, n_6_2684, n_6_2683, 
    n_6_2682, n_6_2681, n_6_2680, n_6_2679, n_6_2678, CLOCK_slo__n58182, n_6_2676, 
    n_6_2675, CLOCK_opt_ipo_n46038, n_6_2673, n_6_2672, slo__sro_n6239, n_6_2670, 
    slo__sro_n15108, n_6_2668, n_6_2667, CLOCK_slo__n56467, n_6_2665}));
datapath__0_132 i_6_31 (.p_2 ({n_6_510, n_6_509, n_6_508, n_6_507, n_6_506, n_6_505, 
    n_6_504, n_6_503, n_6_502, n_6_501, n_6_500, n_6_499, n_6_498, n_6_497, n_6_496, 
    n_6_495, n_6_494, n_6_493, n_6_492, n_6_491, n_6_490, n_6_489, n_6_488, n_6_487, 
    n_6_486, n_6_485, n_6_484, n_6_483, n_6_482, n_6_481, n_6_480, n_6_479}), .p_0 ({
    n_6_30, hfn_ipo_n30, n_6_28, drc_ipo_n26574, n_6_26, n_6_25, CLOCK_sgo__n47054, 
    CLOCK_sgo__n47050, n_6_22, n_6_21, n_6_20, n_6_19, CLOCK_sgo__n47026, n_6_17, 
    n_6_16, n_6_15, n_6_14, n_6_13, n_6_12, n_6_11, n_6_10, drc_ipo_n26591, slo__n26654, 
    slo__n4932, slo__n26805, slo__n26713, slo__n16572, slo__n26761, slo__n3800, slo__n16608, 
    slo__n31700, sgo__n1276}), .p_1 ({uc_14, n_6_2726, n_6_2725, n_6_2724, n_6_2723, 
    n_6_2722, n_6_2721, n_6_2720, slo__n16557, n_6_2718, n_6_2717, n_6_2716, n_6_2715, 
    n_6_2714, n_6_2713, n_6_2712, n_6_2711, n_6_2710, n_6_2709, slo___n16308, n_6_2707, 
    slo___n8747, opt_ipo_n24173, n_6_2704, n_6_2703, n_6_2702, slo__n17720, CLOCK_opt_ipo_n46124, 
    CLOCK_sgo__n47093, n_6_2698, slo__n32451, n_6_2696}), .p_1_3_PP_0 (CLOCK_sgo__n47093));
datapath__0_131 i_6_30 (.p_1 ({n_6_478, n_6_477, n_6_476, n_6_475, n_6_474, n_6_473, 
    n_6_472, n_6_471, n_6_470, n_6_469, n_6_468, n_6_467, n_6_466, n_6_465, n_6_464, 
    n_6_463, n_6_462, n_6_461, n_6_460, n_6_459, n_6_458, n_6_457, n_6_456, n_6_455, 
    n_6_454, n_6_453, n_6_452, n_6_451, n_6_450, n_6_449, n_6_448, n_6_447}), .Multiplier ({
    Multiplier[31], hfn_ipo_n25, Multiplier[29], Multiplier[28], Multiplier[27], 
    drc_ipoPP_6, CLOCK_sgo__n46841, drc_ipo_n26620, drc_ipoPP_5, drc_ipo_n26617, 
    Multiplier[21], Multiplier[20], CLOCK_sgo__n46725, Multiplier[18], drc_ipoPP_4, 
    drc_ipoPP_3, Multiplier[15], drc_ipo_n26609, CLOCK_sgo__n46815, Multiplier[12], 
    Multiplier[11], drc_ipo_n26605, drc_ipoPP_1, drc_ipoPP_0, drc_ipo_n26602, drc_ipo_n26599, 
    drc_ipo_n26600, slo__n4944, slo__n3804, sgo__n1306, drc_ipo_n26598, sgo__n1276})
    , .p_0 ({uc_13, n_6_2726, n_6_2725, n_6_2724, n_6_2723, CLOCK_slo__n55755, n_6_2721, 
    slo__n14626, n_6_2719, slo__n18079, n_6_2717, n_6_2716, n_6_2715, n_6_2714, n_6_2713, 
    n_6_2712, n_6_2711, n_6_2710, n_6_2709, slo__n38783, slo__n38566, slo___n8747, 
    opt_ipo_n24173, slo__n37549, n_6_2703, n_6_2702, n_6_2701, CLOCK_opt_ipo_n46124, 
    CLOCK_sgo__n47093, n_6_2698, slo__n32451, n_6_2696}), .p_0_1_PP_0 (slo__n32451));
datapath__0_127 i_6_27 (.p_2 ({n_6_446, n_6_445, n_6_444, n_6_443, n_6_442, n_6_441, 
    n_6_440, n_6_439, n_6_438, n_6_437, n_6_436, n_6_435, n_6_434, n_6_433, n_6_432, 
    n_6_431, n_6_430, n_6_429, n_6_428, n_6_427, n_6_426, n_6_425, n_6_424, n_6_423, 
    n_6_422, n_6_421, n_6_420, n_6_419, n_6_418, n_6_417, n_6_416, n_6_415}), .p_0 ({
    n_6_30, hfn_ipo_n30, n_6_28, drc_ipo_n26574, n_6_26, n_6_25, CLOCK_sgo__n47054, 
    CLOCK_sgo__n47050, n_6_22, n_6_21, n_6_20, n_6_19, CLOCK_sgo__n47026, n_6_17, 
    n_6_16, n_6_15, n_6_14, n_6_13, n_6_12, n_6_11, n_6_10, drc_ipo_n26591, slo__n26654, 
    slo__n4932, slo__n26805, slo__n26713, slo__n16572, slo__n26761, slo__n3800, slo__n16608, 
    slo__n31700, sgo__n1276}), .p_1 ({uc_12, n_6_2757, n_6_2756, n_6_2755, n_6_2754, 
    opt_ipo_n44116, CLOCK_slo__n56713, n_6_2751, n_6_2750, n_6_2749, n_6_2748, n_6_2747, 
    n_6_2746, slo__n15246, slo__n15241, n_6_2743, n_6_2742, n_6_2741, slo__n15271, 
    n_6_2739, n_6_2738, slo__n18737, slo__n18771, n_6_2735, opt_ipo_n25116, CLOCK_opt_ipo_n45873, 
    n_6_2732, n_6_2731, slo__n15976, slo__n14148, n_6_2728, n_6_2727}));
datapath__0_126 i_6_26 (.p_1 ({n_6_414, n_6_413, n_6_412, n_6_411, n_6_410, n_6_409, 
    n_6_408, n_6_407, n_6_406, n_6_405, n_6_404, n_6_403, n_6_402, n_6_401, n_6_400, 
    n_6_399, n_6_398, n_6_397, n_6_396, n_6_395, n_6_394, n_6_393, n_6_392, n_6_391, 
    n_6_390, n_6_389, n_6_388, n_6_387, n_6_386, n_6_385, n_6_384, n_6_383}), .Multiplier ({
    Multiplier[31], hfn_ipo_n25, Multiplier[29], Multiplier[28], Multiplier[27], 
    drc_ipoPP_6, CLOCK_sgo__n46841, drc_ipo_n26620, drc_ipoPP_5, drc_ipo_n26617, 
    Multiplier[21], Multiplier[20], CLOCK_sgo__n46725, Multiplier[18], drc_ipoPP_4, 
    drc_ipoPP_3, Multiplier[15], drc_ipo_n26609, CLOCK_sgo__n46815, Multiplier[12], 
    Multiplier[11], drc_ipo_n26605, drc_ipoPP_1, drc_ipoPP_0, drc_ipo_n26602, drc_ipo_n26599, 
    drc_ipo_n26600, slo__n4944, slo__n3804, sgo__n1306, drc_ipo_n26598, sgo__n1276})
    , .p_0 ({uc_11, n_6_2757, n_6_2756, n_6_2755, n_6_2754, opt_ipo_n44116, n_6_2752, 
    n_6_2751, slo__n39084, slo__n18877, n_6_2748, n_6_2747, n_6_2746, n_6_2745, n_6_2744, 
    n_6_2743, n_6_2742, n_6_2741, n_6_2740, n_6_2739, n_6_2738, n_6_2737, n_6_2736, 
    n_6_2735, opt_ipo_n25116, CLOCK_opt_ipo_n45873, n_6_2732, n_6_2731, n_6_2730, 
    n_6_2729, n_6_2728, n_6_2727}));
datapath__0_122 i_6_23 (.p_2 ({n_6_382, n_6_381, n_6_380, n_6_379, n_6_378, n_6_377, 
    n_6_376, n_6_375, n_6_374, n_6_373, n_6_372, n_6_371, n_6_370, n_6_369, n_6_368, 
    n_6_367, n_6_366, n_6_365, n_6_364, n_6_363, n_6_362, n_6_361, n_6_360, n_6_359, 
    n_6_358, n_6_357, n_6_356, n_6_355, n_6_354, n_6_353, n_6_352, n_6_351}), .p_0 ({
    n_6_30, hfn_ipo_n30, n_6_28, drc_ipo_n26574, n_6_26, n_6_25, CLOCK_sgo__n47054, 
    CLOCK_sgo__n47050, n_6_22, n_6_21, n_6_20, n_6_19, CLOCK_sgo__n47025, n_6_17, 
    n_6_16, n_6_15, n_6_14, n_6_13, n_6_12, n_6_11, n_6_10, drc_ipo_n26591, slo__n26654, 
    slo__n4932, slo__n26805, slo__n26713, slo__n16572, slo__n26761, slo__n3800, slo__n16608, 
    slo__n31700, sgo__n1276}), .p_1 ({uc_10, n_6_2788, n_6_2787, n_6_2786, n_6_2785, 
    n_6_2784, opt_ipo_n45565, n_6_2782, slo__n16864, n_6_2780, n_6_2779, CLOCK_slo__n56734, 
    n_6_2777, n_6_2776, n_6_2775, n_6_2774, n_6_2773, slo__n18766, slo__n18277, n_6_2770, 
    n_6_2769, slo__n18776, slo__n18465, slo__n18297, slo__sro_n8872, slo__sro_n34940, 
    n_6_2763, CLOCK_slo__n57523, CLOCK_slo__n55377, n_6_2760, CLOCK_slo___n58400, 
    n_6_2758}));
datapath__0_121 i_6_22 (.p_1 ({n_6_350, n_6_349, n_6_348, n_6_347, n_6_346, n_6_345, 
    n_6_344, n_6_343, n_6_342, n_6_341, n_6_340, n_6_339, n_6_338, n_6_337, n_6_336, 
    n_6_335, n_6_334, n_6_333, n_6_332, n_6_331, n_6_330, n_6_329, n_6_328, n_6_327, 
    n_6_326, n_6_325, n_6_324, n_6_323, n_6_322, n_6_321, n_6_320, n_6_319}), .Multiplier ({
    Multiplier[31], hfn_ipo_n25, Multiplier[29], Multiplier[28], Multiplier[27], 
    drc_ipoPP_6, CLOCK_sgo__n46841, drc_ipo_n26620, drc_ipoPP_5, drc_ipo_n26617, 
    Multiplier[21], Multiplier[20], CLOCK_sgo__n46725, Multiplier[18], drc_ipoPP_4, 
    drc_ipoPP_3, Multiplier[15], drc_ipo_n26609, CLOCK_sgo__n46815, Multiplier[12], 
    Multiplier[11], drc_ipo_n26605, drc_ipoPP_1, drc_ipoPP_0, drc_ipo_n26602, drc_ipo_n26599, 
    drc_ipo_n26600, slo__n4944, slo__n3804, sgo__n1306, drc_ipo_n26598, sgo__n1276})
    , .p_0 ({uc_9, CLOCK_slo__n55865, n_6_2787, slo__n16774, slo__n14894, slo__n15162, 
    n_6_1_966, n_6_2782, n_6_2781, n_6_2780, n_6_2779, n_6_2778, n_6_2777, n_6_2776, 
    n_6_2775, n_6_2774, n_6_2773, n_6_2772, n_6_2771, n_6_2770, n_6_2769, n_6_2768, 
    n_6_2767, n_6_2766, slo__sro_n8872, slo__sro_n34940, CLOCK_slo__n57456, n_6_2762, 
    opt_ipo_n24326, n_6_2760, CLOCK_slo___n58400, n_6_2758}), .opt_ipoPP_0 (opt_ipo_n45565));
datapath__0_117 i_6_19 (.p_2 ({n_6_318, n_6_317, n_6_316, n_6_315, n_6_314, n_6_313, 
    n_6_312, n_6_311, n_6_310, n_6_309, n_6_308, n_6_307, n_6_306, n_6_305, n_6_304, 
    n_6_303, n_6_302, n_6_301, n_6_300, n_6_299, n_6_298, n_6_297, n_6_296, n_6_295, 
    n_6_294, n_6_293, n_6_292, n_6_291, n_6_290, n_6_289, n_6_288, n_6_287}), .p_0 ({
    n_6_30, hfn_ipo_n30, n_6_28, drc_ipo_n26574, n_6_26, n_6_25, CLOCK_sgo__n47054, 
    CLOCK_sgo__n47050, n_6_22, n_6_21, n_6_20, n_6_19, CLOCK_sgo__n47025, n_6_17, 
    n_6_16, n_6_15, n_6_14, n_6_13, n_6_12, n_6_11, n_6_10, drc_ipo_n26591, slo__n26654, 
    slo__n4932, slo__n26805, slo__n26713, slo__n16572, slo__n26761, slo__n3800, slo__n16608, 
    slo__n31700, sgo__n1276}), .p_1 ({uc_8, opt_ipo_n25006, n_6_2818, n_6_2817, n_6_2816, 
    n_6_2815, slo___n18581, n_6_2813, n_6_2812, n_6_2811, n_6_2810, slo__n17290, 
    n_6_1_995, n_6_2807, opt_ipo_n24503, n_6_2805, n_6_2804, n_6_2803, n_6_2802, 
    n_6_2801, n_6_2800, n_6_2799, opt_ipo_n25120, n_6_1_984, n_6_2796, n_6_2795, 
    n_6_2794, n_6_2793, n_6_2792, CLOCK_slo__n56313, n_6_2790, CLOCK_slo___n65042}));
datapath__0_116 i_6_18 (.p_1 ({n_6_286, n_6_285, n_6_284, n_6_283, n_6_282, n_6_281, 
    n_6_280, n_6_279, n_6_278, n_6_277, n_6_276, n_6_275, n_6_274, n_6_273, n_6_272, 
    n_6_271, n_6_270, n_6_269, n_6_268, n_6_267, n_6_266, n_6_265, n_6_264, n_6_263, 
    n_6_262, n_6_261, n_6_260, n_6_259, n_6_258, n_6_257, n_6_256, n_6_255}), .Multiplier ({
    Multiplier[31], hfn_ipo_n25, Multiplier[29], Multiplier[28], Multiplier[27], 
    drc_ipoPP_6, CLOCK_sgo__n46841, drc_ipo_n26620, drc_ipoPP_5, drc_ipo_n26617, 
    Multiplier[21], Multiplier[20], CLOCK_sgo__n46725, Multiplier[18], drc_ipoPP_4, 
    drc_ipoPP_3, Multiplier[15], drc_ipo_n26609, drc_ipoPP_2, Multiplier[12], Multiplier[11], 
    drc_ipo_n26605, drc_ipoPP_1, drc_ipoPP_0, drc_ipo_n26602, drc_ipo_n26599, drc_ipo_n26600, 
    slo__n4944, slo__n3804, sgo__n1306, drc_ipo_n26598, sgo__n1276}), .p_0 ({uc_7, 
    opt_ipo_n25007, n_6_2818, slo__n17942, CLOCK_slo__n55860, n_6_2815, slo__n11409, 
    n_6_2813, slo__n15087, n_6_2811, n_6_2810, n_6_2809, n_6_1_995, n_6_2807, opt_ipo_n24503, 
    n_6_2805, n_6_2804, n_6_2803, n_6_2802, n_6_2801, n_6_2800, n_6_2799, opt_ipo_n25120, 
    n_6_1_984, n_6_2796, n_6_2795, n_6_2794, n_6_2793, n_6_2792, CLOCK_slo__n56313, 
    n_6_2790, CLOCK_slo___n65042}), .opt_ipoPP_2 (opt_ipo_n25006));
datapath__0_112 i_6_15 (.p_2 ({n_6_254, n_6_253, n_6_252, n_6_251, n_6_250, n_6_249, 
    n_6_248, n_6_247, n_6_246, n_6_245, n_6_244, n_6_243, n_6_242, n_6_241, n_6_240, 
    n_6_239, n_6_238, n_6_237, n_6_236, n_6_235, n_6_234, n_6_233, n_6_232, n_6_231, 
    n_6_230, n_6_229, n_6_228, n_6_227, n_6_226, n_6_225, n_6_224, n_6_223}), .p_0 ({
    n_6_30, hfn_ipo_n30, n_6_28, drc_ipo_n26574, n_6_26, n_6_25, CLOCK_sgo__n47054, 
    CLOCK_sgo__n47050, n_6_22, n_6_21, n_6_20, n_6_19, CLOCK_sgo__n47025, CLOCK_sgo__n47004, 
    n_6_16, n_6_15, n_6_14, n_6_13, n_6_12, n_6_11, n_6_10, drc_ipo_n26591, slo__n26654, 
    slo__n4932, slo__n26805, slo__n26713, slo__n16572, slo__n26761, slo__n3800, slo__n16608, 
    slo__n31700, sgo__n1276}), .p_1 ({uc_6, n_6_2850, n_6_2849, slo__n18653, slo__n18626, 
    slo__n18732, n_6_2845, n_6_2844, n_6_2843, n_6_2842, slo___n7881, n_6_2840, n_6_2839, 
    CLOCK_slo__n58422, CLOCK_slo___n57806, n_6_2836, n_6_2835, n_6_2834, n_6_2833, 
    n_6_2832, n_6_2831, n_6_2830, n_6_2829, n_6_2828, n_6_2827, n_6_2826, CLOCK_slo__n56284, 
    CLOCK_opt_ipo_n46137, CLOCK_slo__n64837, slo___n5717, n_6_2821, n_6_2820}));
datapath__0_111 i_6_14 (.p_1 ({n_6_222, n_6_221, n_6_220, n_6_219, n_6_218, n_6_217, 
    n_6_216, n_6_215, n_6_214, n_6_213, n_6_212, n_6_211, n_6_210, n_6_209, n_6_208, 
    n_6_207, n_6_206, n_6_205, n_6_204, n_6_203, n_6_202, n_6_201, n_6_200, n_6_199, 
    n_6_198, n_6_197, n_6_196, n_6_195, n_6_194, n_6_193, n_6_192, n_6_191}), .Multiplier ({
    Multiplier[31], hfn_ipo_n25, Multiplier[29], Multiplier[28], Multiplier[27], 
    drc_ipoPP_6, CLOCK_sgo__n46841, drc_ipo_n26620, drc_ipoPP_5, drc_ipo_n26617, 
    Multiplier[21], Multiplier[20], Multiplier[19], Multiplier[18], drc_ipoPP_4, 
    drc_ipoPP_3, Multiplier[15], drc_ipo_n26609, drc_ipoPP_2, Multiplier[12], Multiplier[11], 
    drc_ipo_n26605, drc_ipoPP_1, drc_ipoPP_0, drc_ipo_n26602, drc_ipo_n26599, drc_ipo_n26600, 
    slo__n4944, slo__n3804, sgo__n1306, drc_ipo_n26598, sgo__n1276}), .p_0 ({uc_5, 
    n_6_2850, n_6_2849, n_6_2848, n_6_2847, n_6_2846, n_6_2845, n_6_2844, slo__n14633, 
    n_6_2842, slo___n7881, n_6_2840, n_6_2839, slo___n8281, CLOCK_slo___n57806, n_6_2836, 
    n_6_2835, n_6_2834, n_6_2833, n_6_2832, n_6_2831, n_6_2830, n_6_2829, n_6_2828, 
    n_6_2827, n_6_2826, CLOCK_opt_ipo_n46133, CLOCK_opt_ipo_n46137, opt_ipo_n24190, 
    slo___n5717, n_6_2821, n_6_2820}), .p_0_17_PP_0 (CLOCK_slo___n57806));
datapath__0_107 i_6_11 (.p_2 ({n_6_190, n_6_189, n_6_188, n_6_187, n_6_186, n_6_185, 
    n_6_184, n_6_183, n_6_182, n_6_181, n_6_180, n_6_179, n_6_178, n_6_177, n_6_176, 
    n_6_175, n_6_174, n_6_173, n_6_172, n_6_171, n_6_170, n_6_169, n_6_168, n_6_167, 
    n_6_166, n_6_165, n_6_164, n_6_163, n_6_162, n_6_161, n_6_160, n_6_159}), .p_0 ({
    n_6_30, hfn_ipo_n30, n_6_28, drc_ipo_n26574, n_6_26, n_6_25, CLOCK_sgo__n47054, 
    CLOCK_sgo__n47050, n_6_22, n_6_21, n_6_20, n_6_19, CLOCK_sgo__n47025, CLOCK_sgo__n47004, 
    n_6_16, n_6_15, n_6_14, n_6_13, n_6_12, n_6_11, n_6_10, drc_ipo_n26591, slo__n26654, 
    slo__n4932, slo__n26805, slo__n26713, slo__n16572, slo__n26761, slo__n3800, slo__n16608, 
    slo__n31700, sgo__n1276}), .p_1 ({uc_4, n_6_2881, n_6_2880, n_6_1_1074, slo__sro_n23158, 
    slo__n18727, n_6_2876, slo__n19260, opt_ipo_n24784, slo__n13851, n_6_2872, n_6_2871, 
    slo__n13864, n_6_2869, n_6_2868, n_6_2867, n_6_2866, n_6_2865, n_6_2864, n_6_2863, 
    n_6_2862, n_6_2861, n_6_2860, n_6_2859, n_6_2858, slo__n38665, spw__n68416, n_6_2855, 
    n_6_2854, n_6_2853, n_6_2852, n_6_2851}), .p_0_9_PP_0 (n_6_8));
datapath__0_106 i_6_10 (.p_1 ({n_6_158, n_6_157, n_6_156, n_6_155, n_6_154, n_6_153, 
    n_6_152, n_6_151, n_6_150, n_6_149, n_6_148, n_6_147, n_6_146, n_6_145, n_6_144, 
    n_6_143, n_6_142, n_6_141, n_6_140, n_6_139, n_6_138, n_6_137, n_6_136, n_6_135, 
    n_6_134, n_6_133, n_6_132, n_6_131, n_6_130, n_6_129, n_6_128, n_6_127}), .Multiplier ({
    Multiplier[31], hfn_ipo_n25, Multiplier[29], Multiplier[28], Multiplier[27], 
    drc_ipoPP_6, CLOCK_sgo__n46841, drc_ipo_n26620, drc_ipoPP_5, drc_ipo_n26617, 
    Multiplier[21], Multiplier[20], Multiplier[19], Multiplier[18], drc_ipoPP_4, 
    drc_ipoPP_3, Multiplier[15], drc_ipo_n26609, drc_ipoPP_2, Multiplier[12], Multiplier[11], 
    drc_ipo_n26605, drc_ipoPP_1, drc_ipoPP_0, drc_ipo_n26602, drc_ipo_n26599, drc_ipo_n26600, 
    slo__n4944, slo__n3804, sgo__n1306, drc_ipo_n26598, sgo__n1276}), .p_0 ({uc_3, 
    n_6_2881, n_6_2880, n_6_1_1074, slo__sro_n23158, n_6_2877, n_6_2876, n_6_2875, 
    opt_ipo_n24784, n_6_2873, n_6_2872, n_6_2871, n_6_2870, n_6_2869, n_6_2868, CLOCK_slo__n57483, 
    n_6_2866, n_6_2865, n_6_2864, n_6_2863, n_6_2862, n_6_2861, n_6_2860, CLOCK_slo__n56881, 
    n_6_2858, n_6_2857, spw__n68416, n_6_2855, slo__n10924, slo__sro_n35509, slo__n35483, 
    n_6_2851}));
datapath__0_102 i_6_7 (.p_2 ({n_6_126, n_6_125, n_6_124, n_6_123, n_6_122, n_6_121, 
    n_6_120, n_6_119, n_6_118, n_6_117, n_6_116, n_6_115, n_6_114, n_6_113, n_6_112, 
    n_6_111, n_6_110, n_6_109, n_6_108, n_6_107, n_6_106, n_6_105, n_6_104, n_6_103, 
    n_6_102, n_6_101, n_6_100, n_6_99, n_6_98, n_6_97, n_6_96, n_6_95}), .p_0 ({n_6_30, 
    hfn_ipo_n30, n_6_28, drc_ipo_n26574, n_6_26, n_6_25, CLOCK_sgo__n47054, CLOCK_sgo__n47050, 
    n_6_22, n_6_21, n_6_20, n_6_19, CLOCK_sgo__n47025, CLOCK_sgo__n47003, n_6_16, 
    n_6_15, n_6_14, n_6_13, n_6_12, n_6_11, n_6_10, drc_ipo_n26591, n_6_8, slo__n4932, 
    slo__n26805, slo__n26713, slo__n16572, drc_ipo_n26596, slo__n3800, slo__n38599, 
    drc_ipo_n26597, sgo__n1276}), .p_1 ({uc_2, n_6_2912, n_6_2911, n_6_2910, n_6_2909, 
    n_6_2908, n_6_2907, n_6_2906, n_6_2905, CLOCK_slo__n56075, n_6_2903, slo__n39957, 
    CLOCK_slo__n57534, n_6_2900, n_6_2899, slo__n35792, n_6_2897, n_6_2896, n_6_2895, 
    n_6_2894, n_6_2893, n_6_2892, n_6_2891, n_6_2890, n_6_2889, CLOCK_opt_ipo_n46146, 
    n_6_2887, slo__n36214, slo__n38218, slo__n16550, n_6_2883, CLOCK_spw__n65836})
    , .p_0_9_PP_0 (n_6_8), .opt_ipoPP_2 (opt_ipo_n45480));
datapath__0_101 i_6_6 (.p_1 ({n_6_94, n_6_93, n_6_92, n_6_91, n_6_90, n_6_89, n_6_88, 
    n_6_87, n_6_86, n_6_85, n_6_84, n_6_83, n_6_82, n_6_81, n_6_80, n_6_79, n_6_78, 
    n_6_77, n_6_76, n_6_75, n_6_74, n_6_73, n_6_72, n_6_71, n_6_70, n_6_69, n_6_68, 
    n_6_67, n_6_66, n_6_65, n_6_64, n_6_63}), .Multiplier ({Multiplier[31], hfn_ipo_n25, 
    Multiplier[29], Multiplier[28], Multiplier[27], drc_ipoPP_6, CLOCK_sgo__n46841, 
    drc_ipo_n26620, drc_ipoPP_5, drc_ipo_n26617, Multiplier[21], Multiplier[20], 
    Multiplier[19], Multiplier[18], drc_ipoPP_4, drc_ipoPP_3, Multiplier[15], drc_ipo_n26609, 
    drc_ipoPP_2, Multiplier[12], Multiplier[11], drc_ipo_n26605, drc_ipoPP_1, drc_ipoPP_0, 
    drc_ipo_n26602, drc_ipo_n26599, drc_ipo_n26600, slo__n4944, slo__n3804, sgo__n1306, 
    drc_ipo_n26598, sgo__n1276}), .p_0 ({uc_1, n_6_2912, n_6_2911, n_6_2910, n_6_2909, 
    n_6_2908, n_6_2907, n_6_2906, n_6_2905, n_6_2904, n_6_2903, n_6_2902, n_6_2901, 
    n_6_2900, n_6_2899, n_6_2898, n_6_2897, n_6_2896, n_6_2895, n_6_2894, n_6_2893, 
    n_6_2892, n_6_2891, slo__n12005, n_6_2889, CLOCK_opt_ipo_n46146, n_6_2887, n_6_2886, 
    n_6_2885, n_6_2884, slo__n16791, CLOCK_spw__n65836}), .opt_ipoPP_3 (opt_ipo_n45480));
datapath__0_96 i_6_2 (.p_1 ({n_6_62, n_6_61, n_6_60, n_6_59, n_6_58, n_6_57, n_6_56, 
    n_6_55, n_6_54, n_6_53, n_6_52, n_6_51, n_6_50, n_6_49, n_6_48, n_6_47, n_6_46, 
    n_6_45, n_6_44, n_6_43, n_6_42, n_6_41, n_6_40, n_6_39, n_6_38, n_6_37, n_6_36, 
    n_6_35, n_6_34, n_6_33, n_6_32, n_6_31}), .Multiplier ({Multiplier[31], hfn_ipo_n25, 
    Multiplier[29], Multiplier[28], Multiplier[27], drc_ipoPP_6, CLOCK_sgo__n46841, 
    drc_ipo_n26620, drc_ipoPP_5, drc_ipo_n26617, Multiplier[21], Multiplier[20], 
    Multiplier[19], Multiplier[18], drc_ipoPP_4, drc_ipoPP_3, Multiplier[15], drc_ipo_n26609, 
    drc_ipoPP_2, Multiplier[12], Multiplier[11], drc_ipo_n26605, drc_ipoPP_1, drc_ipoPP_0, 
    drc_ipo_n26602, drc_ipo_n26599, drc_ipo_n26600, slo__n4944, slo__n3804, sgo__n1306, 
    sgo__n1292, sgo__n1276}), .p_0 ({n_6_2913, n_6_30, hfn_ipo_n30, n_6_28, drc_ipo_n26574, 
    n_6_26, n_6_25, CLOCK_sgo__n47054, CLOCK_sgo__n47050, n_6_22, n_6_21, n_6_20, 
    n_6_19, CLOCK_sgo__n47025, CLOCK_sgo__n47003, n_6_16, n_6_15, n_6_14, n_6_13, 
    n_6_12, n_6_11, n_6_10, n_6_9, n_6_8, n_6_7, n_6_6, n_6_5, n_6_4, n_6_3, n_6_2, 
    n_6_1, n_6_0}));
datapath i_6_0 (.p_0 ({n_6_30, n_6_29, n_6_28, n_6_27, n_6_26, n_6_25, n_6_24, CLOCK_sgo__n47050, 
    n_6_22, n_6_21, n_6_20, n_6_19, CLOCK_sgo__n47025, CLOCK_sgo__n47003, n_6_16, 
    n_6_15, n_6_14, n_6_13, n_6_12, n_6_11, n_6_10, n_6_9, n_6_8, n_6_7, n_6_6, n_6_5, 
    n_6_4, n_6_3, n_6_2, n_6_1, n_6_0, uc_0}), .p_0_18_PP_1 (CLOCK_sgo__n47004), .p_0_18_PP_2 (CLOCK_sgo__n47005)
    , .p_0_19_PP_1 (CLOCK_sgo__n47026), .p_0_24_PP_2 (CLOCK_sgo__n47051), .Multiplier ({
    Multiplier[31], hfn_ipo_n26, drc_ipo_n26625, drc_ipo_n26624, drc_ipoPP_7, drc_ipoPP_6, 
    Multiplier[25], drc_ipo_n26620, drc_ipoPP_5, Multiplier[22], drc_ipo_n26616, 
    Multiplier[20], drc_ipo_n26614, drc_ipo_n26613, Multiplier[17], Multiplier[16], 
    drc_ipo_n26610, Multiplier[14], Multiplier[13], Multiplier[12], Multiplier[11], 
    Multiplier[10], drc_ipoPP_1, drc_ipoPP_0, drc_ipo_n26602, Multiplier[6], Multiplier[5], 
    Multiplier[4], Multiplier[3], Multiplier[2], Multiplier[1], Multiplier[0]}), .drc_ipoPP_0 (drc_ipo_n26606));
BUF_X16 hfn_ipo_c25 (.Z (hfn_ipo_n25), .A (Multiplier[30]));
BUF_X16 hfn_ipo_c26 (.Z (hfn_ipo_n26), .A (Multiplier[30]));
BUF_X4 hfn_ipo_c27 (.Z (hfn_ipo_n27), .A (Multiplier[30]));
NAND2_X1 slo__sro_c38983 (.ZN (slo__sro_n35313), .A1 (n_6_1627), .A2 (slo___n23215));
CLKBUF_X3 hfn_ipo_c29 (.Z (hfn_ipo_n29), .A (Multiplier_0_PP_0));
BUF_X16 hfn_ipo_c30 (.Z (hfn_ipo_n30), .A (n_6_29));
BUF_X2 hfn_ipo_c31 (.Z (hfn_ipo_n31), .A (n_6_29));
CLKBUF_X2 hfn_ipo_c32 (.Z (hfn_ipo_n32), .A (n_6_29));
BUF_X16 hfn_ipo_c33 (.Z (hfn_ipo_n33), .A (n_0_0_1));
BUF_X2 hfn_ipo_c34 (.Z (hfn_ipo_n34), .A (n_0_0_1));
BUF_X16 hfn_ipo_c35 (.Z (hfn_ipo_n35), .A (n_0_0_2));
BUF_X2 hfn_ipo_c36 (.Z (hfn_ipo_n36), .A (n_0_0_2));
BUF_X2 sgo__c1051 (.Z (sgo__n1292), .A (slo__n2560));
BUF_X4 sgo__c1077 (.Z (sgo__n1314), .A (n_6_2));
BUF_X32 sgo__c1066 (.Z (sgo__n1306), .A (slo__n2708));
AND2_X1 sgo__sro_c1396 (.ZN (sgo__sro_n1584), .A1 (slo__n30589), .A2 (n_6_4));
AOI21_X1 sgo__sro_c1397 (.ZN (sgo__sro_n1583), .A (sgo__sro_n1584), .B1 (n_6_5), .B2 (opt_ipo_n24358));
BUF_X8 sgo__c1074 (.Z (sgo__n1311), .A (n_6_1));
INV_X1 sgo__sro_c1398 (.ZN (sgo__sro_n1582), .A (sgo__sro_n1583));
AOI21_X2 sgo__sro_c1399 (.ZN (n_6_1_1085), .A (sgo__sro_n1582), .B1 (n_6_36), .B2 (n_6_1_1114));
BUF_X1 sgo__c1027 (.Z (sgo__n1271), .A (n_6_0));
BUF_X16 sgo__c1032 (.Z (sgo__n1276), .A (Multiplier[0]));
NAND2_X1 sgo__sro_c1418 (.ZN (sgo__sro_n1601), .A1 (n_6_3), .A2 (opt_ipo_n24358));
NAND2_X1 sgo__sro_c1419 (.ZN (sgo__sro_n1600), .A1 (sgo__sro_n1602), .A2 (sgo__sro_n1601));
AOI21_X4 sgo__sro_c1420 (.ZN (sgo__sro_n1599), .A (sgo__sro_n1600), .B1 (n_6_34), .B2 (n_6_1_1114));
INV_X1 sgo__sro_c1465 (.ZN (sgo__sro_n1645), .A (opt_ipo_n24358));
NAND2_X1 sgo__sro_c1466 (.ZN (sgo__sro_n1644), .A1 (slo__n4932), .A2 (slo__n30589));
OAI21_X1 sgo__sro_c1467 (.ZN (sgo__sro_n1643), .A (sgo__sro_n1644), .B1 (slo__n26658), .B2 (sgo__sro_n1645));
AOI21_X2 sgo__sro_c1468 (.ZN (n_6_1_1088), .A (sgo__sro_n1643), .B1 (n_6_39), .B2 (n_6_1_1114));
INV_X1 sgo__sro_c1501 (.ZN (sgo__sro_n1676), .A (sgo__sro_n1677));
NAND2_X1 slo__sro_c16813 (.ZN (slo__sro_n15110), .A1 (n_6_2701), .A2 (n_6_1_868));
AOI22_X1 sgo__sro_c1511 (.ZN (sgo__sro_n1688), .A1 (n_6_6), .A2 (opt_ipo_n24358), .B1 (drc_ipo_n26595), .B2 (slo__n30589));
INV_X1 sgo__sro_c1512 (.ZN (sgo__sro_n1687), .A (sgo__sro_n1688));
AOI21_X1 sgo__sro_c1513 (.ZN (sgo__sro_n1686), .A (sgo__sro_n1687), .B1 (n_6_37), .B2 (n_6_1_1114));
AOI21_X1 sgo__sro_c1551 (.ZN (n_6_1_1090), .A (sgo__sro_n1718), .B1 (n_6_41), .B2 (n_6_1_1114));
INV_X1 slo__sro_c2006 (.ZN (slo__sro_n2107), .A (slo__sro_n2108));
AOI21_X4 sgo__sro_c953 (.ZN (sgo__sro_n1215), .A (n_6_1_62), .B1 (n_6_1950), .B2 (n_6_1_64));
INV_X4 sgo__sro_c954 (.ZN (sgo__sro_n1214), .A (sgo__sro_n1215));
AOI21_X2 sgo__sro_c955 (.ZN (sgo__sro_n1213), .A (sgo__sro_n1214), .B1 (n_6_1982), .B2 (n_6_1_65));
INV_X1 slo__sro_c2022 (.ZN (slo__sro_n2122), .A (slo__sro_n2123));
AOI21_X1 slo__sro_c2023 (.ZN (n_6_1_1089), .A (slo__sro_n2122), .B1 (n_6_40), .B2 (n_6_1_1114));
NAND2_X1 slo__sro_c2048 (.ZN (slo__sro_n2144), .A1 (slo__n30589), .A2 (n_6_19));
NAND2_X1 slo__sro_c2049 (.ZN (slo__sro_n2143), .A1 (opt_ipo_n24358), .A2 (n_6_20));
NAND2_X1 slo__sro_c2050 (.ZN (slo__sro_n2142), .A1 (slo__sro_n2144), .A2 (slo__sro_n2143));
AOI22_X4 sgo__sro_c1371 (.ZN (sgo__sro_n1559), .A1 (sgo__n1314), .A2 (sgo__n691), .B1 (sgo__n1311), .B2 (sgo__n711));
NAND2_X1 slo__sro_c41345 (.ZN (slo__sro_n37452), .A1 (slo__sro_n37453), .A2 (slo__sro_n37454));
AOI21_X4 sgo__sro_c1373 (.ZN (sgo__sro_n1557), .A (CLOCK_opt_ipo_n46189), .B1 (n_6_33), .B2 (n_6_1_1114));
INV_X1 slo__sro_c2076 (.ZN (slo__sro_n2165), .A (slo__sro_n2166));
AOI21_X1 slo__sro_c2077 (.ZN (slo__sro_n2164), .A (slo__sro_n2165), .B1 (n_6_43), .B2 (n_6_1_1114));
AOI22_X1 slo__sro_c2107 (.ZN (slo__sro_n2196), .A1 (n_6_11), .A2 (opt_ipo_n24358)
    , .B1 (n_6_10), .B2 (slo__n30589));
INV_X1 slo__sro_c2108 (.ZN (slo__sro_n2195), .A (slo__sro_n2196));
AOI21_X1 slo__sro_c2109 (.ZN (slo__sro_n2194), .A (slo__sro_n2195), .B1 (n_6_42), .B2 (n_6_1_1114));
INV_X1 slo__sro_c2121 (.ZN (slo__sro_n2207), .A (slo__sro_n2208));
AOI21_X1 slo__sro_c2122 (.ZN (slo__sro_n2206), .A (slo__sro_n2207), .B1 (n_6_45), .B2 (n_6_1_1114));
AOI21_X1 slo__sro_c2134 (.ZN (slo__sro_n2221), .A (slo__sro_n2222), .B1 (CLOCK_sgo__n47050), .B2 (opt_ipo_n24358));
INV_X1 slo__sro_c2135 (.ZN (slo__sro_n2220), .A (slo__sro_n2221));
AOI21_X1 slo__sro_c2136 (.ZN (n_6_1_1103), .A (slo__sro_n2220), .B1 (n_6_54), .B2 (n_6_1_1114));
INV_X1 slo__sro_c2148 (.ZN (slo__sro_n2231), .A (slo__sro_n2232));
AOI21_X1 slo__sro_c2149 (.ZN (slo__sro_n2230), .A (slo__sro_n2231), .B1 (n_6_49), .B2 (n_6_1_1114));
NAND2_X1 slo__sro_c2160 (.ZN (slo__sro_n2243), .A1 (n_6_15), .A2 (opt_ipo_n24358));
NAND2_X1 slo__sro_c2161 (.ZN (slo__sro_n2242), .A1 (slo__sro_n2244), .A2 (slo__sro_n2243));
AOI21_X1 slo__sro_c2162 (.ZN (n_6_1_1095), .A (slo__sro_n2242), .B1 (n_6_46), .B2 (n_6_1_1114));
INV_X1 slo__sro_c2174 (.ZN (slo__sro_n2252), .A (slo__sro_n2253));
AOI21_X1 slo__sro_c2175 (.ZN (n_6_1_1097), .A (slo__sro_n2252), .B1 (n_6_48), .B2 (n_6_1_1114));
INV_X1 slo__sro_c2186 (.ZN (slo__sro_n2261), .A (slo__sro_n2262));
AOI21_X1 slo__sro_c2187 (.ZN (slo__sro_n2260), .A (slo__sro_n2261), .B1 (n_6_47), .B2 (n_6_1_1114));
INV_X1 slo__sro_c2198 (.ZN (slo__sro_n2273), .A (slo__sro_n2274));
AOI21_X1 slo__sro_c2199 (.ZN (slo__sro_n2272), .A (slo__sro_n2273), .B1 (n_6_50), .B2 (n_6_1_1114));
NAND2_X1 slo__sro_c2210 (.ZN (slo__sro_n2286), .A1 (opt_ipo_n24358), .A2 (n_6_13));
NAND2_X1 slo__sro_c2211 (.ZN (slo__sro_n2285), .A1 (slo__sro_n2287), .A2 (slo__sro_n2286));
AOI21_X1 slo__sro_c2212 (.ZN (slo__sro_n2284), .A (slo__sro_n2285), .B1 (n_6_44), .B2 (n_6_1_1114));
INV_X1 slo__sro_c2232 (.ZN (slo__sro_n2308), .A (opt_ipo_n24358));
NAND2_X1 slo__sro_c2233 (.ZN (slo__sro_n2307), .A1 (slo__n30589), .A2 (CLOCK_sgo__n47050));
OAI21_X1 slo__sro_c2234 (.ZN (slo__sro_n2306), .A (slo__sro_n2307), .B1 (slo__sro_n2309), .B2 (slo__sro_n2308));
AOI21_X1 slo__sro_c2235 (.ZN (n_6_1_1104), .A (slo__sro_n2306), .B1 (n_6_55), .B2 (n_6_1_1114));
INV_X1 slo__sro_c2248 (.ZN (slo__sro_n2318), .A (slo__sro_n2319));
AOI21_X1 slo__sro_c2249 (.ZN (n_6_1_1102), .A (slo__sro_n2318), .B1 (n_6_53), .B2 (n_6_1_1114));
INV_X1 slo__sro_c2275 (.ZN (slo__sro_n2338), .A (slo__sro_n2339));
AOI21_X1 slo__sro_c2276 (.ZN (n_6_1_1106), .A (slo__sro_n2338), .B1 (n_6_57), .B2 (n_6_1_1114));
INV_X1 slo__sro_c2287 (.ZN (slo__sro_n2347), .A (slo__sro_n2348));
AOI21_X1 slo__sro_c2288 (.ZN (slo__sro_n2346), .A (slo__sro_n2347), .B1 (n_6_52), .B2 (n_6_1_1114));
INV_X2 slo__sro_c2303 (.ZN (slo__sro_n2362), .A (slo__sro_n34792));
AOI21_X4 slo__sro_c2304 (.ZN (n_6_1_1081), .A (slo__sro_n2362), .B1 (n_6_32), .B2 (n_6_1_1114));
INV_X1 slo__sro_c2315 (.ZN (slo__sro_n2371), .A (slo__sro_n2372));
AOI21_X1 slo__sro_c2316 (.ZN (slo__sro_n2370), .A (slo__sro_n2371), .B1 (n_6_58), .B2 (n_6_1_1114));
INV_X1 slo__sro_c2349 (.ZN (slo__sro_n2400), .A (slo__sro_n2401));
AOI21_X1 slo__sro_c2350 (.ZN (n_6_1_1105), .A (slo__sro_n2400), .B1 (n_6_56), .B2 (n_6_1_1114));
INV_X1 slo__sro_c2361 (.ZN (slo__sro_n2409), .A (slo__sro_n2410));
AOI21_X1 slo__sro_c2362 (.ZN (slo__sro_n2408), .A (slo__sro_n2409), .B1 (n_6_59), .B2 (n_6_1_1114));
BUF_X1 slo__c2536 (.Z (slo__n2560), .A (Multiplier[1]));
BUF_X4 slo__c2703 (.Z (slo__n2708), .A (Multiplier[2]));
AOI21_X1 slo__sro_c41346 (.ZN (n_6_1_1004), .A (slo__sro_n37452), .B1 (n_6_252), .B2 (n_6_1_1010));
NAND2_X1 slo__sro_c2996 (.ZN (slo__sro_n2970), .A1 (n_6_2258), .A2 (n_6_1_343));
INV_X1 slo__sro_c2997 (.ZN (slo__sro_n2969), .A (slo__sro_n2970));
AOI21_X1 CLOCK_slo__sro_c69772 (.ZN (n_6_1_951), .A (CLOCK_slo__sro_n62841), .B1 (n_6_266), .B2 (n_6_1_974));
NAND2_X1 slo__sro_c3094 (.ZN (slo__sro_n3058), .A1 (n_6_1_274), .A2 (n_6_1551));
NAND2_X1 slo__sro_c3095 (.ZN (slo__sro_n3057), .A1 (slo__sro_n3058), .A2 (slo__sro_n3059));
AOI21_X2 slo__sro_c3096 (.ZN (slo__sro_n3056), .A (slo__sro_n3057), .B1 (n_6_1583), .B2 (slo___n23244));
BUF_X32 slo__c3926 (.Z (slo__n3800), .A (opt_ipo_n24698));
NAND2_X1 slo__sro_c3871 (.ZN (slo__sro_n3750), .A1 (n_6_1549), .A2 (n_6_1_274));
AOI21_X2 slo__sro_c3873 (.ZN (slo__sro_n3748), .A (slo__sro_n3749), .B1 (n_6_1581), .B2 (slo___n23244));
NAND2_X1 slo__sro_c3872 (.ZN (slo__sro_n3749), .A1 (slo__sro_n3750), .A2 (slo__sro_n3751));
CLKBUF_X2 slo__c3922 (.Z (slo__n3796), .A (n_6_3));
BUF_X32 slo__c3930 (.Z (slo__n3804), .A (Multiplier[3]));
BUF_X4 slo__c3966 (.Z (slo__n3834), .A (n_6_5));
AND2_X1 slo__sro_c4039 (.ZN (slo__sro_n3905), .A1 (n_6_2224), .A2 (n_6_1_308));
NAND2_X1 slo__sro_c3993 (.ZN (slo__sro_n3862), .A1 (n_6_2244), .A2 (n_6_1_343));
INV_X1 CLOCK_slo__sro_c68065 (.ZN (CLOCK_slo__sro_n61296), .A (CLOCK_slo__sro_n61297));
INV_X1 CLOCK_slo__sro_c68077 (.ZN (CLOCK_slo__sro_n61307), .A (CLOCK_slo__sro_n61308));
NAND2_X1 CLOCK_sgo__sro_c51347 (.ZN (CLOCK_sgo__sro_n47134), .A1 (CLOCK_sgo__sro_n47136), .A2 (CLOCK_sgo__sro_n47135));
INV_X1 slo__sro_c4404 (.ZN (slo__sro_n4232), .A (slo__sro_n4233));
AOI221_X2 slo__sro_c4405 (.ZN (n_6_1_682), .A (slo__sro_n4232), .B1 (n_6_789), .B2 (n_6_1_694)
    , .C1 (n_6_821), .C2 (n_6_1_695));
INV_X1 slo__sro_c35179 (.ZN (slo__sro_n31562), .A (slo__sro_n5988));
NAND2_X1 slo__sro_c4465 (.ZN (slo__sro_n4287), .A1 (n_6_1354), .A2 (n_6_1_379));
NAND2_X1 slo__sro_c4466 (.ZN (slo__sro_n4286), .A1 (slo__sro_n4287), .A2 (slo__sro_n4288));
AOI21_X2 slo__sro_c4467 (.ZN (n_6_1_356), .A (slo__sro_n4286), .B1 (n_6_1386), .B2 (n_6_1_380));
NAND2_X1 slo__sro_c4522 (.ZN (slo__sro_n4339), .A1 (slo__sro_n4340), .A2 (slo__sro_n4341));
AOI21_X2 slo__sro_c4523 (.ZN (slo__sro_n4338), .A (slo__sro_n4339), .B1 (n_6_876), .B2 (n_6_1_660));
BUF_X16 sgo__c249 (.Z (n_6_1_695), .A (sgo__n471));
NAND2_X1 slo__sro_c4828 (.ZN (slo__sro_n4616), .A1 (slo__mro_n32529), .A2 (slo__sro_n4618));
AND2_X1 slo__sro_c4494 (.ZN (slo__sro_n4313), .A1 (n_6_2341), .A2 (n_6_1_448));
INV_X1 slo__L1_c1_c43530 (.ZN (slo__n39285), .A (slo__n39286));
AOI21_X1 slo__sro_c4829 (.ZN (slo__sro_n4615), .A (slo__sro_n4616), .B1 (n_6_1768), .B2 (n_6_1_170));
NAND2_X1 slo__sro_c4872 (.ZN (slo__sro_n4661), .A1 (n_6_2166), .A2 (n_6_1_238));
BUF_X16 sgo__c260 (.Z (n_6_1_694), .A (sgo__n482));
BUF_X2 opt_ipo_c49475 (.Z (opt_ipo_n45132), .A (opt_ipo_n45134));
NAND2_X1 slo__sro_c4733 (.ZN (slo__sro_n4530), .A1 (n_6_1_693), .A2 (n_6_2568));
NAND2_X1 slo__sro_c4734 (.ZN (slo__sro_n4529), .A1 (n_6_794), .A2 (n_6_1_694));
NAND2_X1 slo__sro_c4735 (.ZN (slo__sro_n4528), .A1 (slo__sro_n4529), .A2 (slo__sro_n4530));
AOI21_X2 slo__sro_c4736 (.ZN (n_6_1_687), .A (slo__sro_n4528), .B1 (n_6_826), .B2 (n_6_1_695));
AOI222_X1 slo__sro_c39144 (.ZN (slo__sro_n35466), .A1 (n_6_203), .A2 (n_6_1_1009)
    , .B1 (n_6_235), .B2 (n_6_1_1010), .C1 (n_6_2832), .C2 (CLOCK_sgo__n46950));
BUF_X16 sgo__c273 (.Z (n_6_1_730), .A (sgo__n495));
NAND2_X1 slo__sro_c4890 (.ZN (slo__sro_n4672), .A1 (slo__sro_n4673), .A2 (slo__sro_n4674));
AOI21_X1 slo__sro_c4891 (.ZN (n_6_1_1020), .A (slo__sro_n4672), .B1 (n_6_137), .B2 (n_6_1_1044));
AOI21_X4 CLOCK_sgo__sro_c51312 (.ZN (n_6_1_160), .A (CLOCK_sgo__sro_n47109), .B1 (n_6_1784), .B2 (CLOCK_sgo__n48020));
NAND2_X1 slo__sro_c33544 (.ZN (slo__sro_n30020), .A1 (n_6_1_693), .A2 (n_6_2558));
NAND2_X1 slo__sro_c4913 (.ZN (slo__sro_n4691), .A1 (n_6_2163), .A2 (n_6_1_238));
INV_X1 slo__sro_c4914 (.ZN (slo__sro_n4690), .A (slo__sro_n4691));
BUF_X16 sgo__c286 (.Z (n_6_1_729), .A (sgo__n508));
INV_X1 CLOCK_slo__c59668 (.ZN (n_6_1_52), .A (CLOCK_slo__n54298));
INV_X1 slo__sro_c5017 (.ZN (slo__sro_n4786), .A (n_6_1_553));
NOR2_X1 slo__sro_c5018 (.ZN (slo__sro_n4785), .A1 (slo__sro_n4787), .A2 (slo__sro_n4786));
AOI221_X2 slo__sro_c5019 (.ZN (slo__sro_n4784), .A (slo__sro_n4785), .B1 (n_6_1047)
    , .B2 (n_6_1_554), .C1 (n_6_1079), .C2 (slo___n23457));
NAND2_X1 slo__sro_c5047 (.ZN (slo__sro_n4815), .A1 (n_6_1_1080), .A2 (n_6_122));
NAND2_X1 slo__sro_c5048 (.ZN (slo__sro_n4814), .A1 (slo__sro_n4815), .A2 (slo__sro_n4816));
INV_X4 sgo__c299 (.ZN (sgo__n522), .A (sgo__n521));
INV_X16 sgo__c300 (.ZN (n_6_1_765), .A (sgo__n522));
AND2_X2 CLOCK_slo__c70738 (.ZN (CLOCK_slo__sro_n56306), .A1 (n_6_263), .A2 (n_6_1_974));
NAND2_X2 slo__sro_c5085 (.ZN (slo__sro_n4846), .A1 (n_6_1621), .A2 (slo___n23215));
NAND2_X4 slo__sro_c5086 (.ZN (slo__sro_n4845), .A1 (slo__sro_n4846), .A2 (slo__sro_n4847));
AOI21_X1 slo__sro_c5087 (.ZN (slo__sro_n4844), .A (slo__sro_n4845), .B1 (n_6_1653), .B2 (drc_ipo_n26601));
NAND2_X1 slo__sro_c5122 (.ZN (slo__sro_n4882), .A1 (n_6_1137), .A2 (slo___n23268));
NAND2_X1 slo__sro_c5123 (.ZN (slo__sro_n4881), .A1 (slo__sro_n4882), .A2 (slo__sro_n4883));
BUF_X16 sgo__c313 (.Z (n_6_1_764), .A (sgo__n535));
AOI21_X1 slo__sro_c5124 (.ZN (slo__sro_n4880), .A (slo__sro_n4881), .B1 (n_6_1105), .B2 (slo___n23277));
AOI221_X2 CLOCK_slo__sro_c68078 (.ZN (slo__sro_n8949), .A (CLOCK_slo__sro_n61307)
    , .B1 (n_6_162), .B2 (n_6_1_1045), .C1 (n_6_130), .C2 (n_6_1_1044));
BUF_X32 slo__c5189 (.Z (slo__n4944), .A (Multiplier[4]));
AND2_X1 slo__sro_c5263 (.ZN (slo__sro_n5017), .A1 (n_6_2315), .A2 (n_6_1_413));
BUF_X16 sgo__c322 (.Z (n_6_1_800), .A (sgo__n544));
AOI21_X2 CLOCK_slo__sro_c68589 (.ZN (CLOCK_slo__sro_n61783), .A (CLOCK_slo__sro_n61784)
    , .B1 (n_6_1829), .B2 (slo___n23404));
AND2_X1 CLOCK_slo__sro_c52819 (.ZN (CLOCK_slo__sro_n48338), .A1 (n_6_2609), .A2 (n_6_1_763));
BUF_X32 slo__c5199 (.Z (slo__n4958), .A (Multiplier[5]));
NAND2_X1 slo__sro_c5307 (.ZN (slo__sro_n5058), .A1 (n_6_1485), .A2 (n_6_1_309));
BUF_X32 sgo__c331 (.Z (n_6_1_799), .A (sgo__n553));
NAND2_X1 slo__sro_c5308 (.ZN (slo__sro_n5057), .A1 (slo__sro_n5058), .A2 (slo__sro_n5059));
AOI21_X2 slo__sro_c5309 (.ZN (slo__sro_n5056), .A (slo__sro_n5057), .B1 (n_6_1517), .B2 (slo___n23247));
NAND2_X1 CLOCK_slo__sro_c54820 (.ZN (CLOCK_slo__sro_n50131), .A1 (n_6_2460), .A2 (n_6_1_588));
NAND2_X1 slo__sro_c5370 (.ZN (slo__sro_n5119), .A1 (n_6_1_764), .A2 (n_6_658));
NAND2_X1 slo__sro_c5371 (.ZN (slo__sro_n5118), .A1 (slo__sro_n5119), .A2 (slo__sro_n5120));
AOI21_X2 slo__sro_c5372 (.ZN (n_6_1_749), .A (slo__sro_n5118), .B1 (n_6_690), .B2 (n_6_1_765));
BUF_X16 sgo__c344 (.Z (n_6_1_835), .A (sgo__n566));
NAND2_X1 slo__sro_c5490 (.ZN (slo__sro_n5227), .A1 (n_6_1_448), .A2 (n_6_2329));
NAND2_X1 slo__sro_c5491 (.ZN (slo__sro_n5226), .A1 (n_6_1220), .A2 (slo___n23359));
NAND2_X1 slo__sro_c5492 (.ZN (slo__sro_n5225), .A1 (slo__sro_n5226), .A2 (slo__sro_n5227));
INV_X2 slo__c19206 (.ZN (slo__n16984), .A (slo__sro_n20321));
AOI21_X1 CLOCK_slo__sro_c70257 (.ZN (CLOCK_slo__sro_n63268), .A (slo__sro_n11473)
    , .B1 (n_6_303), .B2 (n_6_1_975));
BUF_X16 sgo__c355 (.Z (n_6_1_834), .A (sgo__n577));
NAND2_X1 CLOCK_slo__sro_c56612 (.ZN (CLOCK_slo__sro_n51725), .A1 (n_6_591), .A2 (n_6_1_799));
CLKBUF_X1 spw__L1_c1_c76000 (.Z (CLOCK_slo___n53904), .A (spw__n67799));
INV_X1 CLOCK_slo__sro_c60517 (.ZN (CLOCK_slo__sro_n55022), .A (n_6_1237));
NAND2_X1 slo__sro_c5604 (.ZN (slo__sro_n5333), .A1 (n_6_2584), .A2 (n_6_1_728));
INV_X1 slo__sro_c5605 (.ZN (slo__sro_n5332), .A (slo__sro_n5333));
INV_X1 slo__sro_c20572 (.ZN (slo__sro_n18043), .A (slo__sro_n18044));
INV_X1 slo__sro_c5632 (.ZN (slo__sro_n5353), .A (slo__sro_n5354));
AOI21_X4 CLOCK_slo__sro_c66387 (.ZN (CLOCK_slo__sro_n59842), .A (CLOCK_slo__sro_n59843)
    , .B1 (n_6_871), .B2 (n_6_1_660));
BUF_X16 sgo__c372 (.Z (n_6_1_870), .A (sgo__n594));
NAND2_X1 CLOCK_sgo__sro_c51663 (.ZN (CLOCK_sgo__sro_n47395), .A1 (n_6_738), .A2 (n_6_1_730));
BUF_X32 drc_ipo_c29959 (.Z (drc_ipo_n26582), .A (CLOCK_sgo__n47025));
INV_X1 slo__sro_c36146 (.ZN (slo__sro_n32473), .A (slo__sro_n20127));
INV_X1 slo__sro_c24028 (.ZN (slo__sro_n20923), .A (slo__sro_n20924));
INV_X1 slo__sro_c6033 (.ZN (slo__sro_n5712), .A (n_6_1_553));
NOR2_X1 slo__sro_c6034 (.ZN (slo__sro_n5711), .A1 (slo__sro_n5713), .A2 (slo__sro_n5712));
BUF_X16 sgo__c385 (.Z (n_6_1_869), .A (sgo__n607));
AND2_X1 CLOCK_slo__sro_c59418 (.ZN (CLOCK_slo__sro_n54099), .A1 (CLOCK_slo__sro_n54100), .A2 (CLOCK_slo__sro_n54101));
BUF_X16 sgo__c388 (.Z (n_6_1_905), .A (sgo__n610));
NAND2_X1 slo__sro_c6219 (.ZN (slo__sro_n5877), .A1 (slo___n23215), .A2 (n_6_1609));
BUF_X16 sgo__c391 (.Z (n_6_1_904), .A (sgo__n613));
NAND2_X1 slo__sro_c41070 (.ZN (slo__sro_n37209), .A1 (slo__sro_n37210), .A2 (slo__sro_n37211));
AND2_X1 slo__sro_c6186 (.ZN (slo__sro_n5844), .A1 (n_6_2403), .A2 (n_6_1_518));
BUF_X16 sgo__c396 (.Z (n_6_1_940), .A (sgo__n618));
NAND2_X1 slo__sro_c6220 (.ZN (slo__sro_n5876), .A1 (slo__sro_n5877), .A2 (slo__sro_n5878));
BUF_X16 sgo__c399 (.Z (n_6_1_939), .A (sgo__n621));
AOI222_X2 slo__sro_c6134 (.ZN (slo__sro_n5794), .A1 (n_6_1133), .A2 (slo___n23268)
    , .B1 (n_6_1101), .B2 (slo___n23277), .C1 (slo___n15030), .C2 (n_6_1_518));
AOI221_X2 slo__sro_c6254 (.ZN (slo__sro_n5907), .A (slo__sro_n5908), .B1 (n_6_1676)
    , .B2 (slo___n23239), .C1 (n_6_1708), .C2 (slo___n23407));
NAND2_X1 slo__sro_c6313 (.ZN (slo__sro_n5964), .A1 (n_6_682), .A2 (n_6_1_765));
NAND2_X1 slo__sro_c6314 (.ZN (slo__sro_n5963), .A1 (slo__sro_n5964), .A2 (slo__sro_n5965));
BUF_X16 sgo__c408 (.Z (n_6_1_975), .A (sgo__n630));
AND2_X1 slo__sro_c6294 (.ZN (slo__sro_n5946), .A1 (n_6_2268), .A2 (n_6_1_378));
NAND2_X1 CLOCK_sgo__sro_c51787 (.ZN (CLOCK_sgo__sro_n47501), .A1 (CLOCK_sgo__sro_n47502), .A2 (CLOCK_sgo__sro_n47503));
INV_X1 slo__sro_c35287 (.ZN (slo__sro_n31656), .A (CLOCK_sgo__n46945));
BUF_X16 sgo__c415 (.Z (n_6_1_974), .A (sgo__n637));
INV_X1 slo__sro_c23913 (.ZN (slo__sro_n20820), .A (n_6_2653));
NAND2_X1 slo__sro_c6398 (.ZN (slo__sro_n6041), .A1 (n_6_2330), .A2 (n_6_1_448));
INV_X4 sgo__c422 (.ZN (sgo__n645), .A (sgo__n644));
INV_X16 sgo__c423 (.ZN (n_6_1_1010), .A (sgo__n645));
NAND2_X1 slo__sro_c6399 (.ZN (slo__sro_n6040), .A1 (n_6_1221), .A2 (slo___n23359));
NAND2_X1 slo__sro_c40224 (.ZN (slo__sro_n36477), .A1 (slo__sro_n36478), .A2 (slo__sro_n36479));
AOI21_X2 slo__sro_c6401 (.ZN (slo__sro_n6038), .A (slo__sro_n6039), .B1 (n_6_1253), .B2 (slo___n23274));
NAND2_X2 slo__sro_c6530 (.ZN (slo__sro_n6162), .A1 (n_6_1_309), .A2 (n_6_1478));
NAND2_X2 slo__sro_c6531 (.ZN (slo__sro_n6161), .A1 (slo__sro_n6162), .A2 (slo__sro_n6163));
BUF_X16 sgo__c434 (.Z (n_6_1_1009), .A (sgo__n656));
AOI21_X4 slo__sro_c6532 (.ZN (slo__sro_n6160), .A (slo__sro_n6161), .B1 (n_6_1510), .B2 (slo___n23247));
BUF_X16 sgo__c437 (.Z (n_6_1_1045), .A (sgo__n659));
NAND2_X1 slo__sro_c6612 (.ZN (slo__sro_n6241), .A1 (n_6_454), .A2 (n_6_1_869));
NAND2_X1 slo__sro_c6560 (.ZN (slo__sro_n6194), .A1 (n_6_2301), .A2 (n_6_1_413));
NAND2_X1 slo__sro_c6561 (.ZN (slo__sro_n6193), .A1 (n_6_1287), .A2 (n_6_1_414));
BUF_X16 sgo__c444 (.Z (n_6_1_1044), .A (sgo__n666));
NAND2_X1 slo__sro_c6562 (.ZN (slo__sro_n6192), .A1 (slo__sro_n6193), .A2 (slo__sro_n6194));
AOI21_X2 slo__sro_c6563 (.ZN (slo__sro_n6191), .A (slo__sro_n6192), .B1 (n_6_1319), .B2 (slo___n43257));
AOI21_X2 slo__sro_c6614 (.ZN (CLOCK_slo__n48618), .A (slo__sro_n6240), .B1 (n_6_486), .B2 (n_6_1_870));
NAND2_X1 CLOCK_slo__sro_c71926 (.ZN (CLOCK_slo__sro_n64639), .A1 (n_6_2023), .A2 (n_6_1_98));
INV_X8 sgo__c453 (.ZN (sgo__n676), .A (sgo__n675));
INV_X32 sgo__c454 (.ZN (n_6_1_1080), .A (sgo__n676));
INV_X1 slo__sro_c6744 (.ZN (slo__sro_n6370), .A (n_6_1804));
INV_X1 slo__sro_c6745 (.ZN (slo__sro_n6369), .A (n_6_1_134));
AND2_X1 slo__sro_c6660 (.ZN (slo__sro_n6283), .A1 (n_6_2346), .A2 (n_6_1_448));
NAND2_X1 CLOCK_slo__sro_c60594 (.ZN (CLOCK_slo__sro_n55086), .A1 (slo___n23229), .A2 (n_6_1412));
OAI21_X1 slo__sro_c6747 (.ZN (slo__sro_n6367), .A (slo__sro_n6368), .B1 (slo__sro_n6370), .B2 (slo__sro_n6369));
INV_X8 sgo__c465 (.ZN (sgo__n688), .A (sgo__n687));
INV_X32 sgo__c466 (.ZN (n_6_1_1079), .A (sgo__n688));
AOI21_X2 slo__sro_c6748 (.ZN (slo__sro_n6366), .A (slo__sro_n6367), .B1 (n_6_1836), .B2 (n_6_1_135));
NOR2_X2 CLOCK_slo__sro_c63592 (.ZN (slo__sro_n8450), .A1 (CLOCK_slo__sro_n57490), .A2 (slo__sro_n8451));
INV_X1 slo__sro_c35470 (.ZN (slo__sro_n31831), .A (slo__sro_n31832));
NAND2_X1 slo__sro_c6915 (.ZN (slo__sro_n6521), .A1 (n_6_118), .A2 (n_6_1_1080));
NAND2_X1 slo__sro_c6916 (.ZN (slo__sro_n6520), .A1 (slo__sro_n6521), .A2 (slo__sro_n6522));
AOI21_X1 slo__sro_c6917 (.ZN (slo__sro_n6519), .A (slo__sro_n6520), .B1 (n_6_86), .B2 (n_6_1_1079));
AOI21_X2 slo__sro_c7050 (.ZN (slo__sro_n6653), .A (slo__sro_n6654), .B1 (n_6_1286), .B2 (n_6_1_414));
NAND2_X1 slo__sro_c6898 (.ZN (slo__sro_n6506), .A1 (n_6_2350), .A2 (n_6_1_448));
NAND2_X2 slo__sro_c6899 (.ZN (slo__sro_n6505), .A1 (n_6_1241), .A2 (slo___n23359));
NAND2_X2 slo__sro_c6900 (.ZN (slo__sro_n6504), .A1 (slo__sro_n6505), .A2 (slo__sro_n6506));
NAND2_X1 slo__sro_c6843 (.ZN (slo__sro_n6457), .A1 (n_6_2136), .A2 (n_6_1_203));
NAND2_X2 slo__sro_c6844 (.ZN (slo__sro_n6456), .A1 (n_6_1692), .A2 (n_6_1_204));
BUF_X32 drc_ipo_c29953 (.Z (drc_ipo_n26576), .A (n_6_22));
NAND2_X2 slo__sro_c6845 (.ZN (slo__sro_n6455), .A1 (slo__sro_n6456), .A2 (slo__sro_n6457));
INV_X1 sgo__c492 (.ZN (sgo__n715), .A (sgo__n714));
INV_X16 sgo__c493 (.ZN (n_6_1_1114), .A (sgo__n715));
AOI21_X2 slo__sro_c6846 (.ZN (n_6_1_199), .A (slo__sro_n6455), .B1 (n_6_1724), .B2 (slo___n23407));
NAND2_X1 slo__sro_c6975 (.ZN (slo__sro_n6578), .A1 (n_6_1667), .A2 (n_6_1_204));
NAND2_X1 slo__sro_c6976 (.ZN (slo__sro_n6577), .A1 (slo__sro_n6578), .A2 (slo__sro_n6579));
NAND2_X1 CLOCK_slo__sro_c67497 (.ZN (CLOCK_slo__sro_n60778), .A1 (n_6_1_168), .A2 (slo__sro_n30921));
INV_X1 slo__sro_c7033 (.ZN (slo__sro_n6638), .A (n_6_2237));
INV_X1 slo__sro_c7034 (.ZN (slo__sro_n6637), .A (n_6_1_343));
NOR2_X1 slo__sro_c7035 (.ZN (slo__sro_n6636), .A1 (slo__sro_n6638), .A2 (slo__sro_n6637));
INV_X1 slo__sro_c45432 (.ZN (slo__sro_n40962), .A (n_6_2637));
NAND2_X2 slo__sro_c7076 (.ZN (slo__sro_n6675), .A1 (n_6_1282), .A2 (n_6_1_414));
NAND2_X2 slo__sro_c7077 (.ZN (slo__sro_n6674), .A1 (slo__sro_n6675), .A2 (slo__sro_n6676));
AOI21_X4 slo__sro_c7078 (.ZN (slo__sro_n6673), .A (slo__sro_n6674), .B1 (n_6_1314), .B2 (slo___n43257));
NAND2_X1 slo__sro_c7092 (.ZN (slo__sro_n6690), .A1 (n_6_1283), .A2 (n_6_1_414));
NAND2_X1 slo__sro_c7093 (.ZN (slo__sro_n6689), .A1 (slo__sro_n6690), .A2 (slo__sro_n6691));
AND2_X1 CLOCK_slo__sro_c60133 (.ZN (CLOCK_slo__sro_n54698), .A1 (n_6_316), .A2 (n_6_1_975));
AND2_X1 slo__sro_c7212 (.ZN (slo__sro_n6791), .A1 (n_6_2308), .A2 (n_6_1_413));
NAND2_X1 slo__sro_c7116 (.ZN (slo__sro_n6708), .A1 (n_6_2429), .A2 (n_6_1_553));
INV_X1 slo__sro_c7117 (.ZN (slo__sro_n6707), .A (slo__sro_n6708));
AOI221_X2 slo__sro_c7118 (.ZN (n_6_1_532), .A (slo__sro_n6707), .B1 (n_6_1035), .B2 (n_6_1_554)
    , .C1 (n_6_1067), .C2 (slo___n23457));
AND2_X2 slo__sro_c44253 (.ZN (slo__sro_n39872), .A1 (n_6_1468), .A2 (n_6_1_345));
AOI21_X2 slo__sro_c7252 (.ZN (slo__sro_n6827), .A (slo__sro_n6828), .B1 (n_6_1228), .B2 (slo___n23359));
NAND2_X1 slo__sro_c7184 (.ZN (slo__sro_n6765), .A1 (n_6_1_343), .A2 (n_6_2247));
NAND2_X1 slo__sro_c7185 (.ZN (slo__sro_n6764), .A1 (slo___n23229), .A2 (n_6_1423));
NAND2_X1 slo__sro_c7186 (.ZN (slo__sro_n6763), .A1 (slo__sro_n6764), .A2 (slo__sro_n6765));
NAND2_X1 CLOCK_slo__sro_c66262 (.ZN (CLOCK_slo__sro_n59730), .A1 (opt_ipo_n45107), .A2 (n_6_1_98));
AOI222_X2 slo__sro_c7274 (.ZN (slo__sro_n6852), .A1 (n_6_1028), .A2 (slo___n23353)
    , .B1 (n_6_1060), .B2 (slo___n23457), .C1 (n_6_2422), .C2 (n_6_1_553));
NAND2_X1 slo__sro_c7293 (.ZN (slo__sro_n6870), .A1 (slo__sro_n6871), .A2 (slo__sro_n6872));
AOI21_X2 slo__sro_c7294 (.ZN (slo__sro_n6869), .A (slo__sro_n6870), .B1 (n_6_1204), .B2 (slo___n23466));
AND2_X1 CLOCK_slo__sro_c54772 (.ZN (CLOCK_slo__sro_n50083), .A1 (n_6_2243), .A2 (n_6_1_343));
AOI21_X1 CLOCK_slo__sro_c72472 (.ZN (CLOCK_slo__sro_n65088), .A (CLOCK_slo__sro_n65089)
    , .B1 (n_6_204), .B2 (n_6_1_1009));
BUF_X8 drc_ipo_c29974 (.Z (drc_ipo_n26597), .A (slo__n5306));
NAND2_X1 slo__sro_c34642 (.ZN (slo__sro_n31052), .A1 (n_6_1298), .A2 (n_6_1_414));
NAND2_X1 CLOCK_slo__sro_c55891 (.ZN (CLOCK_slo__sro_n51095), .A1 (opt_ipo_n24166), .A2 (n_6_1_763));
NAND2_X1 slo__sro_c7517 (.ZN (slo__sro_n7075), .A1 (n_6_1_273), .A2 (n_6_2196));
AOI221_X2 slo__sro_c35289 (.ZN (slo__sro_n31654), .A (slo__sro_n31655), .B1 (n_6_163)
    , .B2 (n_6_1_1045), .C1 (n_6_131), .C2 (n_6_1_1044));
NAND2_X1 slo__sro_c7519 (.ZN (slo__sro_n7073), .A1 (slo__mro_n31601), .A2 (slo__sro_n7075));
AOI21_X2 slo__sro_c7520 (.ZN (n_6_1_267), .A (slo__sro_n7073), .B1 (n_6_1594), .B2 (slo___n23244));
AOI222_X2 slo__sro_c7387 (.ZN (slo__sro_n6955), .A1 (n_6_449), .A2 (n_6_1_869), .B1 (n_6_481)
    , .B2 (n_6_1_870), .C1 (n_6_2698), .C2 (n_6_1_868));
NAND2_X2 slo__sro_c7657 (.ZN (slo__sro_n7188), .A1 (n_6_995), .A2 (slo___n23218));
NAND2_X1 slo__sro_c7461 (.ZN (slo__sro_n7020), .A1 (n_6_2507), .A2 (n_6_1_623));
NAND2_X1 slo__sro_c7462 (.ZN (slo__sro_n7019), .A1 (n_6_923), .A2 (slo___n23367));
NAND2_X1 slo__sro_c7463 (.ZN (slo__sro_n7018), .A1 (slo__sro_n7019), .A2 (slo__sro_n7020));
AOI21_X2 slo__sro_c7464 (.ZN (slo__sro_n7017), .A (slo__sro_n7018), .B1 (n_6_955), .B2 (n_6_1_625));
AOI21_X2 slo__sro_c7659 (.ZN (slo__sro_n7186), .A (slo__sro_n7187), .B1 (n_6_963), .B2 (slo___n23232));
NAND2_X1 slo__sro_c7801 (.ZN (slo__sro_n7334), .A1 (slo__n35802), .A2 (n_6_1_553));
NAND2_X1 slo__sro_c7802 (.ZN (slo__sro_n7333), .A1 (n_6_1033), .A2 (slo___n23353));
AOI222_X2 slo__sro_c7871 (.ZN (slo__sro_n7395), .A1 (n_6_781), .A2 (n_6_1_694), .B1 (n_6_813)
    , .B2 (n_6_1_695), .C1 (n_6_2555), .C2 (n_6_1_693));
NAND2_X1 slo__sro_c7882 (.ZN (slo__sro_n7407), .A1 (n_6_1034), .A2 (slo___n23353));
AOI222_X2 slo__sro_c7689 (.ZN (slo__sro_n7219), .A1 (n_6_525), .A2 (n_6_1_834), .B1 (n_6_557)
    , .B2 (n_6_1_835), .C1 (n_6_2679), .C2 (CLOCK_sgo__n46922));
AOI222_X2 slo__sro_c7631 (.ZN (n_6_1_522), .A1 (n_6_1025), .A2 (slo___n23353), .B1 (n_6_1057)
    , .B2 (slo___n23457), .C1 (n_6_2419), .C2 (n_6_1_553));
INV_X1 CLOCK_sgo__sro_c51363 (.ZN (CLOCK_sgo__sro_n47150), .A (slo__sro_n34361));
NAND2_X1 slo__sro_c7803 (.ZN (slo__sro_n7332), .A1 (slo__sro_n7333), .A2 (slo__sro_n7334));
AOI21_X2 slo__sro_c7804 (.ZN (slo__sro_n7331), .A (slo__sro_n7332), .B1 (n_6_1065), .B2 (slo___n23457));
AOI21_X2 slo__sro_c7884 (.ZN (CLOCK_slo__n55041), .A (slo__sro_n7406), .B1 (n_6_1066), .B2 (slo___n23457));
INV_X1 slo__sro_c7898 (.ZN (slo__sro_n7422), .A (slo__sro_n7423));
NAND2_X1 CLOCK_slo__sro_c65308 (.ZN (CLOCK_slo__sro_n58846), .A1 (CLOCK_slo__sro_n58847), .A2 (CLOCK_slo__sro_n50682));
NAND2_X1 slo__sro_c7777 (.ZN (slo__sro_n7308), .A1 (n_6_1361), .A2 (n_6_1_379));
NAND2_X1 slo__sro_c7778 (.ZN (slo__sro_n7307), .A1 (slo__sro_n7308), .A2 (slo__sro_n7309));
NAND2_X1 slo__sro_c23984 (.ZN (slo__sro_n20888), .A1 (n_6_2508), .A2 (n_6_1_623));
NAND2_X1 slo__sro_c7944 (.ZN (slo__sro_n7467), .A1 (n_6_1_483), .A2 (n_6_2359));
NAND2_X1 slo__sro_c7945 (.ZN (slo__sro_n7466), .A1 (n_6_1155), .A2 (slo___n23364));
AOI21_X1 slo__sro_c7947 (.ZN (n_6_1_454), .A (slo__sro_n7465), .B1 (n_6_1187), .B2 (slo___n23466));
NAND2_X1 slo__sro_c41384 (.ZN (slo__sro_n37484), .A1 (n_6_494), .A2 (n_6_1_870));
AOI222_X2 slo__sro_c8133 (.ZN (slo__sro_n7633), .A1 (n_6_1062), .A2 (slo___n23457)
    , .B1 (n_6_1030), .B2 (slo___n23353), .C1 (n_6_2424), .C2 (n_6_1_553));
AOI21_X1 slo__sro_c8202 (.ZN (slo__sro_n7689), .A (slo__sro_n7690), .B1 (n_6_1006), .B2 (slo___n23218));
NAND2_X1 slo__sro_c8291 (.ZN (slo__sro_n7775), .A1 (CLOCK_opt_ipo_n46133), .A2 (CLOCK_sgo__n46950));
INV_X1 slo__c8272 (.ZN (slo__n7753), .A (n_6_1_791));
NAND2_X2 slo__sro_c8200 (.ZN (slo__sro_n7691), .A1 (n_6_974), .A2 (slo___n23232));
NAND2_X2 CLOCK_slo__sro_c54349 (.ZN (CLOCK_slo__sro_n49713), .A1 (n_6_1193), .A2 (slo___n23466));
AOI222_X2 slo__sro_c8001 (.ZN (slo__sro_n7515), .A1 (n_6_857), .A2 (slo___n23463)
    , .B1 (n_6_889), .B2 (slo___n23451), .C1 (slo___n9717), .C2 (n_6_1_658));
NAND2_X1 slo__sro_c8293 (.ZN (slo__sro_n7773), .A1 (slo__sro_n7774), .A2 (slo__sro_n7775));
AOI21_X1 slo__sro_c8294 (.ZN (slo__sro_n7772), .A (slo__sro_n7773), .B1 (n_6_196), .B2 (n_6_1_1009));
AOI222_X2 slo__sro_c8047 (.ZN (slo__sro_n7557), .A1 (n_6_842), .A2 (slo___n23463)
    , .B1 (n_6_874), .B2 (n_6_1_660), .C1 (opt_ipo_n23804), .C2 (n_6_1_658));
AOI222_X2 slo__sro_c8037 (.ZN (n_6_1_825), .A1 (n_6_568), .A2 (n_6_1_835), .B1 (n_6_536)
    , .B2 (n_6_1_834), .C1 (n_6_2690), .C2 (CLOCK_sgo__n46922));
NAND2_X1 CLOCK_slo__sro_c54348 (.ZN (CLOCK_slo__sro_n49714), .A1 (n_6_2365), .A2 (n_6_1_483));
NAND2_X1 slo__sro_c8353 (.ZN (slo__sro_n7833), .A1 (slo__sro_n7834), .A2 (slo__sro_n7835));
BUF_X8 slo___L1_c26574 (.Z (slo___n23215), .A (n_6_1_239));
NAND2_X1 slo__sro_c8439 (.ZN (slo__sro_n7912), .A1 (n_6_1_799), .A2 (n_6_596));
AND2_X1 slo__sro_c22433 (.ZN (slo__sro_n19450), .A1 (n_6_2565), .A2 (n_6_1_693));
BUF_X4 drc_ipo_c29962 (.Z (drc_ipo_n26585), .A (n_6_16));
AND2_X1 slo__sro_c8426 (.ZN (slo__sro_n7899), .A1 (n_6_2704), .A2 (n_6_1_868));
AOI221_X2 slo__sro_c8427 (.ZN (slo__sro_n7898), .A (slo__sro_n7899), .B1 (n_6_455)
    , .B2 (n_6_1_869), .C1 (n_6_487), .C2 (n_6_1_870));
AND2_X1 slo__sro_c8460 (.ZN (slo__sro_n7933), .A1 (n_6_2763), .A2 (CLOCK_sgo__n46937));
NAND2_X1 CLOCK_sgo__sro_c51533 (.ZN (CLOCK_sgo__sro_n47287), .A1 (n_6_1353), .A2 (n_6_1_379));
NAND2_X1 slo__sro_c8474 (.ZN (slo__sro_n7945), .A1 (slo__sro_n7946), .A2 (slo__sro_n7947));
INV_X2 CLOCK_slo__c60448 (.ZN (CLOCK_slo__n54964), .A (slo__sro_n5855));
INV_X1 slo__sro_c8489 (.ZN (slo__sro_n7960), .A (slo__sro_n7961));
AOI221_X2 slo__sro_c8490 (.ZN (n_6_1_754), .A (slo__sro_n7960), .B1 (n_6_663), .B2 (n_6_1_764)
    , .C1 (n_6_695), .C2 (n_6_1_765));
NAND2_X1 slo__sro_c8570 (.ZN (slo__sro_n8030), .A1 (n_6_2597), .A2 (n_6_1_728));
NAND2_X1 slo__sro_c8571 (.ZN (slo__sro_n8029), .A1 (n_6_728), .A2 (n_6_1_729));
NAND2_X1 slo__sro_c8572 (.ZN (slo__sro_n8028), .A1 (slo__sro_n8029), .A2 (slo__sro_n8030));
AOI21_X1 slo__sro_c8573 (.ZN (n_6_1_720), .A (slo__sro_n8028), .B1 (n_6_760), .B2 (n_6_1_730));
INV_X1 slo__sro_c8593 (.ZN (slo__sro_n8046), .A (slo__sro_n8047));
AOI221_X2 slo__sro_c8594 (.ZN (n_6_1_744), .A (slo__sro_n8046), .B1 (n_6_685), .B2 (n_6_1_765)
    , .C1 (n_6_653), .C2 (n_6_1_764));
AOI222_X2 slo__sro_c8642 (.ZN (slo__sro_n8092), .A1 (n_6_1046), .A2 (n_6_1_554), .B1 (n_6_1078)
    , .B2 (slo___n23457), .C1 (CLOCK_slo__n53562), .C2 (n_6_1_553));
NAND2_X1 CLOCK_slo__sro_c72469 (.ZN (CLOCK_slo__sro_n65091), .A1 (CLOCK_sgo__n46950), .A2 (n_6_2833));
BUF_X4 drc_ipo_c29964 (.Z (drc_ipo_n26587), .A (n_6_13));
AOI221_X2 CLOCK_slo__sro_c69953 (.ZN (CLOCK_slo__sro_n63004), .A (CLOCK_slo__sro_n63005)
    , .B1 (n_6_1041), .B2 (n_6_1_554), .C1 (n_6_1073), .C2 (slo___n23457));
NAND2_X1 slo__sro_c8867 (.ZN (slo__sro_n8297), .A1 (slo__n14626), .A2 (n_6_1_868));
NAND2_X1 slo__sro_c8868 (.ZN (slo__sro_n8296), .A1 (n_6_471), .A2 (n_6_1_869));
NAND2_X1 slo__sro_c8869 (.ZN (slo__sro_n8295), .A1 (slo__sro_n8296), .A2 (slo__sro_n8297));
AOI222_X2 slo__sro_c8803 (.ZN (n_6_1_788), .A1 (n_6_630), .A2 (n_6_1_800), .B1 (n_6_598)
    , .B2 (n_6_1_799), .C1 (n_6_2657), .C2 (n_6_1_798));
INV_X1 slo__sro_c8884 (.ZN (slo__sro_n8310), .A (slo__sro_n8311));
AOI221_X2 slo__sro_c8885 (.ZN (slo__n29454), .A (slo__sro_n8310), .B1 (n_6_666), .B2 (n_6_1_764)
    , .C1 (n_6_698), .C2 (n_6_1_765));
NAND2_X1 slo__sro_c8918 (.ZN (slo__sro_n8340), .A1 (slo__n13799), .A2 (n_6_2906));
NAND2_X1 slo__sro_c8919 (.ZN (slo__sro_n8339), .A1 (n_6_119), .A2 (n_6_1_1080));
AOI21_X1 slo__sro_c8921 (.ZN (n_6_1_1069), .A (slo__sro_n8338), .B1 (n_6_87), .B2 (n_6_1_1079));
NAND2_X1 slo__sro_c8941 (.ZN (slo__sro_n8357), .A1 (n_6_115), .A2 (n_6_1_1080));
NAND2_X1 slo__sro_c8942 (.ZN (slo__sro_n8356), .A1 (slo__sro_n8357), .A2 (slo__sro_n8358));
INV_X1 slo__sro_c44293 (.ZN (slo__sro_n39899), .A (slo__sro_n39900));
NAND2_X1 slo__sro_c8957 (.ZN (slo__sro_n8369), .A1 (n_6_1_1080), .A2 (n_6_117));
NAND2_X1 slo__sro_c8958 (.ZN (slo__sro_n8368), .A1 (slo__sro_n8369), .A2 (slo__sro_n8370));
AOI21_X2 slo__sro_c8959 (.ZN (n_6_1_1067), .A (slo__sro_n8368), .B1 (n_6_85), .B2 (n_6_1_1079));
NAND2_X1 slo__sro_c8983 (.ZN (slo__sro_n8391), .A1 (n_6_70), .A2 (n_6_1_1079));
NAND2_X1 slo__sro_c8984 (.ZN (slo__sro_n8390), .A1 (slo__sro_n8391), .A2 (slo__sro_n8392));
AOI21_X2 slo__sro_c8985 (.ZN (n_6_1_1052), .A (slo__sro_n8390), .B1 (n_6_102), .B2 (n_6_1_1080));
NAND2_X1 slo__sro_c8999 (.ZN (slo__sro_n8403), .A1 (n_6_1_1080), .A2 (n_6_116));
NAND2_X1 slo__sro_c9000 (.ZN (slo__sro_n8402), .A1 (slo__sro_n8403), .A2 (slo__sro_n8404));
AOI21_X1 slo__sro_c9001 (.ZN (n_6_1_1066), .A (slo__sro_n8402), .B1 (n_6_84), .B2 (n_6_1_1079));
NAND2_X1 slo__sro_c9015 (.ZN (slo__sro_n8416), .A1 (n_6_1_1080), .A2 (n_6_114));
NAND2_X1 slo__sro_c9016 (.ZN (slo__sro_n8415), .A1 (slo__sro_n8416), .A2 (slo__sro_n8417));
INV_X1 slo__sro_c44413 (.ZN (slo__sro_n40010), .A (slo__sro_n6636));
NAND2_X1 slo__sro_c9031 (.ZN (slo__sro_n8431), .A1 (n_6_1_1080), .A2 (n_6_121));
NAND2_X2 slo__sro_c9032 (.ZN (slo__sro_n8430), .A1 (slo__sro_n8431), .A2 (slo__sro_n8432));
NAND2_X1 CLOCK_slo__sro_c61708 (.ZN (CLOCK_slo__sro_n56019), .A1 (n_6_2873), .A2 (CLOCK_sgo__n46945));
NAND2_X1 slo__sro_c9055 (.ZN (slo__sro_n8452), .A1 (n_6_1_1080), .A2 (n_6_113));
NAND2_X1 slo__sro_c9056 (.ZN (slo__sro_n8451), .A1 (slo__sro_n8452), .A2 (slo__sro_n8453));
NAND2_X1 CLOCK_slo__sro_c63883 (.ZN (CLOCK_slo__sro_n57701), .A1 (n_6_1_274), .A2 (n_6_1566));
NAND2_X1 slo__sro_c9195 (.ZN (slo__sro_n8581), .A1 (n_6_1_1080), .A2 (n_6_112));
NAND2_X1 slo__sro_c9196 (.ZN (slo__sro_n8580), .A1 (slo__sro_n8581), .A2 (slo__sro_n8582));
AND2_X1 slo__sro_c9095 (.ZN (slo__sro_n8489), .A1 (n_6_2715), .A2 (n_6_1_868));
AOI221_X2 slo__sro_c9096 (.ZN (slo__sro_n8488), .A (slo__sro_n8489), .B1 (n_6_498)
    , .B2 (n_6_1_870), .C1 (n_6_466), .C2 (n_6_1_869));
NAND2_X1 CLOCK_slo__sro_c53149 (.ZN (CLOCK_slo__sro_n48635), .A1 (CLOCK_slo__sro_n48636), .A2 (slo__sro_n18492));
AOI21_X2 CLOCK_slo__sro_c53150 (.ZN (CLOCK_slo__sro_n48634), .A (CLOCK_slo__sro_n48635)
    , .B1 (n_6_453), .B2 (n_6_1_869));
AOI21_X1 slo__sro_c9223 (.ZN (slo__sro_n8602), .A (slo__sro_n8603), .B1 (n_6_66), .B2 (n_6_1_1079));
NAND2_X2 CLOCK_sgo__sro_c51311 (.ZN (CLOCK_sgo__sro_n47109), .A1 (CLOCK_sgo__sro_n47110), .A2 (CLOCK_sgo__sro_n47111));
AOI222_X2 slo__sro_c38958 (.ZN (slo__sro_n35288), .A1 (n_6_308), .A2 (n_6_1_975), .B1 (n_6_276)
    , .B2 (n_6_1_974), .C1 (n_6_2810), .C2 (n_6_1_973));
AOI222_X2 slo__sro_c9275 (.ZN (slo__sro_n8646), .A1 (n_6_822), .A2 (n_6_1_695), .B1 (n_6_790)
    , .B2 (n_6_1_694), .C1 (n_6_2564), .C2 (n_6_1_693));
NAND2_X1 slo__sro_c9323 (.ZN (slo__sro_n8684), .A1 (slo__sro_n8685), .A2 (slo__sro_n8686));
AOI21_X1 slo__sro_c9324 (.ZN (n_6_1_593), .A (slo__sro_n8684), .B1 (n_6_898), .B2 (slo___n23367));
NAND2_X1 slo__sro_c9434 (.ZN (slo__sro_n8778), .A1 (n_6_2862), .A2 (CLOCK_sgo__n46945));
NAND2_X1 slo__sro_c9435 (.ZN (slo__sro_n8777), .A1 (n_6_1_1045), .A2 (n_6_170));
NAND2_X2 CLOCK_slo__sro_c53510 (.ZN (CLOCK_slo__sro_n48958), .A1 (CLOCK_slo__sro_n48959), .A2 (CLOCK_slo__sro_n48960));
AOI222_X2 slo__sro_c9356 (.ZN (n_6_1_648), .A1 (n_6_854), .A2 (slo___n23463), .B1 (n_6_886)
    , .B2 (slo___n23451), .C1 (n_6_2533), .C2 (n_6_1_658));
NAND2_X1 slo__sro_c9419 (.ZN (slo__sro_n8765), .A1 (n_6_530), .A2 (n_6_1_834));
NAND2_X1 slo__sro_c9420 (.ZN (slo__sro_n8764), .A1 (slo__sro_n8765), .A2 (slo__sro_n8766));
NAND2_X1 CLOCK_slo__sro_c62809 (.ZN (CLOCK_slo__sro_n56895), .A1 (n_6_1673), .A2 (slo___n23239));
INV_X1 slo__sro_c30989 (.ZN (slo__sro_n27584), .A (slo__sro_n8057));
NAND2_X1 slo__sro_c9583 (.ZN (slo__sro_n8918), .A1 (n_6_803), .A2 (n_6_1_695));
NAND2_X1 slo__sro_c9538 (.ZN (slo__sro_n8875), .A1 (n_6_1_984), .A2 (n_6_1_973));
NAND2_X1 slo__sro_c9539 (.ZN (slo__sro_n8874), .A1 (n_6_1_975), .A2 (n_6_295));
NAND2_X1 slo__sro_c9540 (.ZN (slo__sro_n8873), .A1 (slo__sro_n8874), .A2 (slo__sro_n8875));
NAND2_X1 CLOCK_slo__sro_c62146 (.ZN (CLOCK_slo__sro_n56378), .A1 (n_6_1_834), .A2 (n_6_534));
NAND2_X1 slo__sro_c9567 (.ZN (slo__sro_n8902), .A1 (n_6_1167), .A2 (slo___n23364));
NAND2_X1 slo__sro_c9568 (.ZN (slo__sro_n8901), .A1 (slo__sro_n8902), .A2 (slo__sro_n8903));
AOI21_X2 slo__sro_c9569 (.ZN (slo__sro_n8900), .A (slo__sro_n8901), .B1 (n_6_1199), .B2 (slo___n23466));
AOI21_X1 slo__sro_c9585 (.ZN (slo__sro_n8916), .A (slo__sro_n8917), .B1 (n_6_771), .B2 (n_6_1_694));
AND2_X1 slo__sro_c9631 (.ZN (slo__sro_n8966), .A1 (opt_ipo_n44116), .A2 (CLOCK_sgo__n46934));
NAND2_X1 slo__sro_c37455 (.ZN (slo__sro_n33778), .A1 (n_6_2476), .A2 (n_6_1_588));
NOR2_X2 CLOCK_slo__sro_c67484 (.ZN (CLOCK_slo__sro_n60762), .A1 (slo__sro_n6577), .A2 (CLOCK_slo__sro_n60763));
NAND2_X1 slo__sro_c9658 (.ZN (slo__sro_n8993), .A1 (n_6_1_1079), .A2 (n_6_69));
NAND2_X1 slo__sro_c9659 (.ZN (slo__sro_n8992), .A1 (slo__sro_n8993), .A2 (slo__sro_n8994));
AOI21_X2 slo__sro_c9660 (.ZN (slo__sro_n8991), .A (slo__sro_n8992), .B1 (n_6_101), .B2 (n_6_1_1080));
NAND2_X1 slo__sro_c9674 (.ZN (slo__sro_n9009), .A1 (n_6_99), .A2 (n_6_1_1080));
NAND2_X2 slo__sro_c9675 (.ZN (slo__sro_n9008), .A1 (slo__sro_n9009), .A2 (slo__sro_n9010));
AOI21_X2 slo__sro_c9676 (.ZN (slo__sro_n9007), .A (slo__sro_n9008), .B1 (n_6_67), .B2 (n_6_1_1079));
NAND2_X1 slo__sro_c9695 (.ZN (slo__sro_n9030), .A1 (n_6_2768), .A2 (CLOCK_sgo__n46937));
INV_X1 slo__sro_c9696 (.ZN (slo__sro_n9029), .A (slo__sro_n9030));
AOI221_X2 slo__sro_c9697 (.ZN (n_6_1_915), .A (slo__sro_n9029), .B1 (n_6_361), .B2 (n_6_1_940)
    , .C1 (n_6_329), .C2 (n_6_1_939));
AOI222_X2 slo__sro_c9748 (.ZN (slo__sro_n9075), .A1 (n_6_869), .A2 (n_6_1_660), .B1 (n_6_837)
    , .B2 (slo___n23463), .C1 (slo___n6972), .C2 (n_6_1_658));
NAND2_X1 slo__sro_c9796 (.ZN (slo__sro_n9123), .A1 (n_6_1359), .A2 (n_6_1_379));
NAND2_X1 slo__sro_c9797 (.ZN (slo__sro_n9122), .A1 (slo__sro_n9123), .A2 (slo__sro_n9124));
AOI21_X2 slo__sro_c9798 (.ZN (n_6_1_361), .A (slo__sro_n9122), .B1 (n_6_1391), .B2 (n_6_1_380));
NAND2_X1 slo__sro_c9874 (.ZN (slo__sro_n9197), .A1 (n_6_2254), .A2 (n_6_1_343));
NAND2_X1 slo__sro_c9875 (.ZN (slo__sro_n9196), .A1 (n_6_1430), .A2 (slo___n23229));
NAND2_X1 slo__sro_c9876 (.ZN (slo__sro_n9195), .A1 (slo__sro_n9196), .A2 (slo__sro_n9197));
AOI21_X2 slo__sro_c9877 (.ZN (slo__sro_n9194), .A (slo__sro_n9195), .B1 (n_6_1462), .B2 (n_6_1_345));
NAND2_X1 slo__sro_c9926 (.ZN (slo__sro_n9244), .A1 (n_6_1284), .A2 (n_6_1_414));
NAND2_X1 slo__sro_c9927 (.ZN (slo__sro_n9243), .A1 (slo__sro_n9244), .A2 (slo__sro_n9245));
AOI21_X2 slo__sro_c9928 (.ZN (slo__sro_n9242), .A (slo__sro_n9243), .B1 (n_6_1316), .B2 (slo___n43257));
AOI221_X2 slo__sro_c10033 (.ZN (slo__sro_n9341), .A (slo__sro_n9342), .B1 (n_6_362)
    , .B2 (n_6_1_940), .C1 (n_6_330), .C2 (n_6_1_939));
AOI21_X4 slo__sro_c46340 (.ZN (slo__sro_n41830), .A (slo__sro_n41831), .B1 (n_6_219), .B2 (n_6_1_1009));
AND2_X1 slo__sro_c10082 (.ZN (slo__sro_n9390), .A1 (n_6_1_238), .A2 (n_6_2142));
NAND2_X1 slo__sro_c23101 (.ZN (slo__sro_n20068), .A1 (CLOCK_sgo__n46937), .A2 (n_6_2782));
NAND2_X1 slo__sro_c35302 (.ZN (slo__sro_n31672), .A1 (n_6_2818), .A2 (n_6_1_973));
NAND2_X1 slo__sro_c10172 (.ZN (slo__sro_n9470), .A1 (n_6_1668), .A2 (slo___n23239));
NAND2_X1 slo__sro_c10173 (.ZN (slo__sro_n9469), .A1 (slo__sro_n9470), .A2 (slo__sro_n9471));
NAND2_X1 CLOCK_slo__sro_c53263 (.ZN (CLOCK_slo__sro_n48742), .A1 (n_6_2146), .A2 (n_6_1_238));
AOI221_X2 slo__sro_c10238 (.ZN (slo__sro_n9533), .A (slo__sro_n9534), .B1 (n_6_1370)
    , .B2 (n_6_1_379), .C1 (n_6_1402), .C2 (n_6_1_380));
INV_X2 slo__L1_c2_c30809 (.ZN (slo__n27410), .A (slo__n27411));
NAND2_X1 slo__sro_c10381 (.ZN (slo__sro_n9672), .A1 (n_6_293), .A2 (n_6_1_975));
NAND2_X1 slo__sro_c10382 (.ZN (slo__sro_n9671), .A1 (slo__sro_n9672), .A2 (slo__sro_n9673));
AOI21_X2 slo__sro_c10383 (.ZN (n_6_1_946), .A (slo__sro_n9671), .B1 (n_6_261), .B2 (n_6_1_974));
AOI21_X2 CLOCK_slo__sro_c56941 (.ZN (CLOCK_slo__sro_n51979), .A (CLOCK_slo__sro_n51980)
    , .B1 (n_6_1136), .B2 (slo___n23268));
NAND2_X2 slo__sro_c10485 (.ZN (slo__sro_n9755), .A1 (n_6_1431), .A2 (slo___n23229));
NAND2_X1 slo__sro_c10433 (.ZN (slo__sro_n9711), .A1 (slo__sro_n9712), .A2 (slo__sro_n9713));
AOI21_X2 slo__sro_c10434 (.ZN (n_6_1_945), .A (slo__sro_n9711), .B1 (n_6_260), .B2 (n_6_1_974));
NAND2_X1 slo__sro_c10484 (.ZN (slo__sro_n9756), .A1 (n_6_2255), .A2 (n_6_1_343));
NAND2_X2 slo__sro_c10486 (.ZN (slo__sro_n9754), .A1 (slo__sro_n9755), .A2 (slo__sro_n9756));
AND2_X1 slo__sro_c10472 (.ZN (slo__sro_n9745), .A1 (n_6_2467), .A2 (n_6_1_588));
AND2_X1 slo__sro_c40748 (.ZN (slo__sro_n36933), .A1 (n_6_2710), .A2 (n_6_1_868));
NAND2_X1 slo__sro_c10528 (.ZN (slo__sro_n9794), .A1 (n_6_2260), .A2 (n_6_1_343));
NOR2_X2 CLOCK_slo__sro_c56214 (.ZN (CLOCK_slo__sro_n51387), .A1 (CLOCK_slo__sro_n51388), .A2 (slo__sro_n16001));
NAND2_X1 CLOCK_slo__sro_c56309 (.ZN (CLOCK_slo__sro_n51474), .A1 (n_6_1694), .A2 (n_6_1_204));
AND2_X1 slo__sro_c44282 (.ZN (slo__sro_n39889), .A1 (n_6_83), .A2 (n_6_1_1079));
NAND2_X1 CLOCK_slo__sro_c58031 (.ZN (CLOCK_slo__sro_n52916), .A1 (slo___n23430), .A2 (n_6_1758));
NAND2_X1 slo__sro_c10617 (.ZN (slo__sro_n9875), .A1 (n_6_2532), .A2 (n_6_1_658));
NAND2_X1 slo__sro_c10618 (.ZN (slo__sro_n9874), .A1 (n_6_885), .A2 (slo___n23451));
NAND2_X1 slo__sro_c10619 (.ZN (slo__sro_n9873), .A1 (slo__sro_n9874), .A2 (slo__sro_n9875));
OAI21_X2 slo__mro_c36700 (.ZN (slo__mro_n33030), .A (slo__sro_n7708), .B1 (slo__mro_n33032), .B2 (slo__mro_n33031));
NAND2_X1 slo__sro_c10730 (.ZN (slo__sro_n9978), .A1 (n_6_1048), .A2 (n_6_1_554));
NAND2_X1 slo__sro_c10731 (.ZN (slo__sro_n9977), .A1 (slo__sro_n9978), .A2 (slo__sro_n9979));
AOI21_X2 slo__sro_c10732 (.ZN (n_6_1_545), .A (slo__sro_n9977), .B1 (n_6_1080), .B2 (slo___n23457));
AND2_X1 slo__sro_c32878 (.ZN (slo__sro_n29381), .A1 (n_6_2215), .A2 (n_6_1_308));
AOI222_X2 slo__sro_c10754 (.ZN (n_6_1_718), .A1 (n_6_726), .A2 (n_6_1_729), .B1 (n_6_758)
    , .B2 (n_6_1_730), .C1 (n_6_2595), .C2 (n_6_1_728));
AOI221_X2 slo__sro_c31253 (.ZN (slo__sro_n27836), .A (slo__sro_n27837), .B1 (n_6_291)
    , .B2 (n_6_1_975), .C1 (n_6_259), .C2 (n_6_1_974));
INV_X1 slo__sro_c10870 (.ZN (slo__sro_n10099), .A (CLOCK_sgo__n46934));
NOR2_X1 slo__sro_c10871 (.ZN (slo__sro_n10098), .A1 (slo__sro_n10100), .A2 (slo__sro_n10099));
INV_X1 slo__sro_c38259 (.ZN (slo__sro_n34623), .A (n_6_2562));
INV_X1 slo__c10950 (.ZN (slo__n10168), .A (n_6_1_760));
AND2_X1 slo__sro_c33208 (.ZN (slo__sro_n29693), .A1 (n_6_2866), .A2 (CLOCK_sgo__n46945));
AOI21_X2 slo__sro_c11069 (.ZN (slo__sro_n10270), .A (slo__sro_n10271), .B1 (n_6_586), .B2 (n_6_1_799));
AND2_X1 CLOCK_slo__sro_c61735 (.ZN (CLOCK_slo__sro_n56037), .A1 (n_6_508), .A2 (n_6_1_870));
INV_X1 slo__c11133 (.ZN (slo__n10331), .A (n_6_1_489));
AOI222_X1 slo__sro_c11110 (.ZN (slo__sro_n10311), .A1 (n_6_1802), .A2 (n_6_1_134)
    , .B1 (n_6_1834), .B2 (n_6_1_135), .C1 (n_6_2056), .C2 (n_6_1_133));
BUF_X1 slo__L2_c3_c34249 (.Z (slo__n30670), .A (slo__n30671));
AOI222_X2 slo__sro_c10990 (.ZN (n_6_1_950), .A1 (n_6_297), .A2 (n_6_1_975), .B1 (n_6_265)
    , .B2 (n_6_1_974), .C1 (n_6_2799), .C2 (n_6_1_973));
NAND2_X1 slo__sro_c11256 (.ZN (slo__sro_n10428), .A1 (n_6_1307), .A2 (n_6_1_414));
AOI21_X2 slo__sro_c11258 (.ZN (slo__sro_n10426), .A (slo__sro_n10427), .B1 (n_6_1339), .B2 (slo___n43257));
AOI221_X2 slo__sro_c11291 (.ZN (n_6_1_442), .A (slo__sro_n10458), .B1 (n_6_1242), .B2 (slo___n23359)
    , .C1 (n_6_1274), .C2 (slo___n23274));
AND2_X1 slo__sro_c37978 (.ZN (slo__sro_n34361), .A1 (n_6_2576), .A2 (n_6_1_728));
AND2_X1 slo__sro_c11178 (.ZN (slo__sro_n10370), .A1 (n_6_2662), .A2 (n_6_1_798));
INV_X1 CLOCK_slo__sro_c56120 (.ZN (CLOCK_slo__sro_n51309), .A (slo__sro_n29693));
NAND2_X2 slo__sro_c33167 (.ZN (slo__sro_n29652), .A1 (n_6_1285), .A2 (n_6_1_414));
NAND2_X2 slo__sro_c11417 (.ZN (slo__sro_n10560), .A1 (slo__sro_n10562), .A2 (slo__sro_n10561));
AOI21_X2 slo__sro_c11418 (.ZN (n_6_1_127), .A (slo__sro_n10560), .B1 (n_6_1850), .B2 (n_6_1_135));
NAND2_X1 slo__sro_c11528 (.ZN (slo__sro_n10651), .A1 (n_6_1819), .A2 (slo___n23226));
NAND2_X1 slo__sro_c35979 (.ZN (slo__sro_n32319), .A1 (n_6_2176), .A2 (n_6_1_273));
NAND2_X1 slo__sro_c11574 (.ZN (slo__sro_n10694), .A1 (n_6_2055), .A2 (n_6_1_133));
NAND2_X1 slo__sro_c11552 (.ZN (slo__sro_n10676), .A1 (n_6_2070), .A2 (n_6_1_133));
NAND2_X1 slo__sro_c11553 (.ZN (slo__sro_n10675), .A1 (n_6_1816), .A2 (n_6_1_134));
NAND2_X1 slo__sro_c11554 (.ZN (slo__sro_n10674), .A1 (slo__sro_n10675), .A2 (slo__sro_n10676));
AOI21_X2 slo__sro_c11555 (.ZN (n_6_1_125), .A (slo__sro_n10674), .B1 (n_6_1848), .B2 (n_6_1_135));
INV_X1 slo__c11512 (.ZN (slo__n10634), .A (n_6_1_139));
AND2_X1 CLOCK_slo__sro_c67483 (.ZN (CLOCK_slo__sro_n60763), .A1 (n_6_1699), .A2 (slo___n23407));
NAND2_X1 CLOCK_sgo__sro_c52005 (.ZN (CLOCK_sgo__sro_n47683), .A1 (CLOCK_opt_ipo_n45779), .A2 (n_6_1_273));
NAND2_X1 slo__sro_c11662 (.ZN (slo__sro_n10770), .A1 (slo__sro_n10772), .A2 (slo__sro_n10771));
INV_X1 slo__c11619 (.ZN (slo__n10734), .A (n_6_1_70));
AOI21_X2 slo__sro_c11663 (.ZN (slo__sro_n10769), .A (slo__sro_n10770), .B1 (n_6_1849), .B2 (n_6_1_135));
AOI222_X2 slo__sro_c11682 (.ZN (n_6_1_824), .A1 (n_6_535), .A2 (n_6_1_834), .B1 (n_6_567)
    , .B2 (n_6_1_835), .C1 (n_6_2689), .C2 (CLOCK_sgo__n46922));
NAND2_X1 CLOCK_slo__sro_c68076 (.ZN (CLOCK_slo__sro_n61308), .A1 (n_6_2854), .A2 (CLOCK_sgo__n46945));
AOI21_X4 CLOCK_slo__sro_c54308 (.ZN (CLOCK_slo__sro_n49672), .A (CLOCK_slo__sro_n49673)
    , .B1 (n_6_1380), .B2 (n_6_1_380));
INV_X1 slo__c11816 (.ZN (slo__n10924), .A (slo__n14340));
INV_X1 slo__c11824 (.ZN (slo__n10929), .A (slo__sro_n6651));
NAND2_X1 slo__sro_c12063 (.ZN (slo__sro_n11125), .A1 (n_6_1157), .A2 (slo___n23364));
AND2_X1 slo__sro_c11851 (.ZN (slo__sro_n10956), .A1 (opt_ipo_n45565), .A2 (CLOCK_sgo__n46937));
BUF_X4 slo__c46252 (.Z (n_6_1_554), .A (slo__n41748));
AND2_X1 slo__sro_c11793 (.ZN (slo__sro_n10905), .A1 (n_6_2802), .A2 (n_6_1_973));
AOI221_X2 CLOCK_slo__sro_c54773 (.ZN (CLOCK_slo__sro_n50082), .A (CLOCK_slo__sro_n50083)
    , .B1 (n_6_1419), .B2 (slo___n23229), .C1 (n_6_1451), .C2 (n_6_1_345));
AND2_X1 slo__sro_c11945 (.ZN (slo__sro_n11035), .A1 (n_6_2803), .A2 (n_6_1_973));
AOI21_X2 CLOCK_sgo__sro_c52082 (.ZN (n_6_1_281), .A (CLOCK_sgo__sro_n47732), .B1 (n_6_1509), .B2 (slo___n23247));
NAND2_X1 slo__sro_c33832 (.ZN (slo__sro_n30287), .A1 (n_6_2398), .A2 (n_6_1_518));
INV_X2 CLOCK_opt_ipo_c50087 (.ZN (CLOCK_opt_ipo_n45744), .A (n_6_1_115));
AOI221_X2 CLOCK_slo__sro_c71382 (.ZN (CLOCK_slo__sro_n64180), .A (CLOCK_slo__sro_n59303)
    , .B1 (n_6_1324), .B2 (slo___n43257), .C1 (n_6_1292), .C2 (n_6_1_414));
NAND2_X1 slo__sro_c12169 (.ZN (slo__sro_n11218), .A1 (CLOCK_sgo__n46922), .A2 (opt_ipo_n44105));
AOI21_X4 slo__mro_c36920 (.ZN (slo__mro_n33266), .A (slo__mro_n33269), .B1 (slo__mro_n33268), .B2 (slo__mro_n33267));
NAND2_X2 slo__mro_c36954 (.ZN (slo__mro_n33301), .A1 (n_6_1980), .A2 (n_6_1_65));
AOI21_X2 slo__sro_c12172 (.ZN (slo__sro_n11215), .A (slo__sro_n11216), .B1 (n_6_569), .B2 (n_6_1_835));
NAND2_X1 slo__sro_c12301 (.ZN (slo__sro_n11319), .A1 (CLOCK_sgo__n46945), .A2 (n_6_2864));
NAND2_X1 slo__sro_c12302 (.ZN (slo__sro_n11318), .A1 (n_6_140), .A2 (n_6_1_1044));
INV_X1 slo__c12115 (.ZN (slo__n11164), .A (CLOCK_slo__sro_n50657));
NAND2_X1 slo__sro_c12303 (.ZN (slo__sro_n11317), .A1 (slo__sro_n11318), .A2 (slo__sro_n11319));
INV_X2 slo__c12248 (.ZN (slo__n11270), .A (n_6_1_789));
AOI21_X2 slo__sro_c12304 (.ZN (n_6_1_1023), .A (slo__sro_n11317), .B1 (n_6_172), .B2 (n_6_1_1045));
INV_X1 slo__c12429 (.ZN (slo__n11420), .A (slo__sro_n28419));
INV_X1 slo__c12439 (.ZN (slo__n11427), .A (slo__sro_n7617));
NAND2_X1 slo__sro_c12450 (.ZN (slo__sro_n11436), .A1 (slo__sro_n11437), .A2 (slo__sro_n11438));
AOI21_X2 slo__sro_c12451 (.ZN (n_6_1_492), .A (slo__sro_n11436), .B1 (n_6_1094), .B2 (slo___n23277));
NAND2_X1 slo__sro_c12489 (.ZN (slo__sro_n11474), .A1 (n_6_2805), .A2 (n_6_1_973));
INV_X1 slo__sro_c41283 (.ZN (slo__sro_n37405), .A (slo__sro_n7478));
NAND2_X2 CLOCK_slo__mro_c70606 (.ZN (CLOCK_slo__mro_n63532), .A1 (n_6_1331), .A2 (slo___n43257));
INV_X1 slo__c12514 (.ZN (slo__n11487), .A (n_6_1_394));
NAND2_X1 slo__sro_c12764 (.ZN (slo__sro_n11709), .A1 (n_6_2863), .A2 (CLOCK_sgo__n46945));
NAND2_X1 slo__sro_c12637 (.ZN (slo__sro_n11595), .A1 (slo__sro_n11596), .A2 (slo__sro_n11597));
AOI21_X2 slo__sro_c12638 (.ZN (slo__sro_n11594), .A (slo__sro_n11595), .B1 (n_6_1340), .B2 (slo___n43257));
AOI221_X2 slo__sro_c12687 (.ZN (n_6_1_513), .A (slo__sro_n11641), .B1 (n_6_1115), .B2 (slo___n23277)
    , .C1 (n_6_1147), .C2 (slo___n23268));
INV_X2 slo__c12225 (.ZN (slo__n11253), .A (slo__sro_n16910));
INV_X2 slo__c13664 (.ZN (slo__n12473), .A (n_6_1_861));
INV_X2 slo__c12726 (.ZN (slo__n11671), .A (n_6_1_295));
NAND2_X1 slo__sro_c12766 (.ZN (slo__sro_n11707), .A1 (slo__sro_n11708), .A2 (slo__sro_n11709));
AND2_X1 slo__sro_c12674 (.ZN (slo__sro_n11633), .A1 (n_6_2444), .A2 (n_6_1_553));
AOI221_X2 slo__sro_c12675 (.ZN (n_6_1_547), .A (slo__sro_n11633), .B1 (n_6_1050), .B2 (n_6_1_554)
    , .C1 (n_6_1082), .C2 (slo___n23457));
AND2_X1 slo__sro_c12786 (.ZN (slo__sro_n11729), .A1 (opt_ipo_n45324), .A2 (n_6_1_203));
AOI221_X2 slo__sro_c12787 (.ZN (slo__sro_n11728), .A (slo__sro_n11729), .B1 (n_6_1717)
    , .B2 (slo___n23407), .C1 (n_6_1685), .C2 (n_6_1_204));
AND2_X1 slo__sro_c12807 (.ZN (slo__sro_n11746), .A1 (n_6_2779), .A2 (CLOCK_sgo__n46937));
AOI221_X2 slo__sro_c12808 (.ZN (n_6_1_926), .A (slo__sro_n11746), .B1 (n_6_372), .B2 (n_6_1_940)
    , .C1 (n_6_340), .C2 (n_6_1_939));
NAND2_X1 slo__sro_c12867 (.ZN (slo__sro_n11797), .A1 (slo__sro_n11798), .A2 (slo__sro_n11799));
INV_X1 slo__sro_c12849 (.ZN (slo__sro_n11786), .A (slo___n18581));
INV_X1 slo__sro_c12850 (.ZN (slo__sro_n11785), .A (n_6_1_973));
NOR2_X1 slo__sro_c12851 (.ZN (slo__sro_n11784), .A1 (slo__sro_n11786), .A2 (slo__sro_n11785));
NAND2_X1 slo__sro_c26177 (.ZN (slo__sro_n22875), .A1 (CLOCK_sgo__n46945), .A2 (n_6_2868));
NAND2_X1 slo__sro_c12897 (.ZN (slo__sro_n11831), .A1 (n_6_2781), .A2 (CLOCK_sgo__n46937));
NAND2_X2 slo__sro_c12898 (.ZN (slo__sro_n11830), .A1 (n_6_342), .A2 (n_6_1_939));
NAND2_X2 slo__sro_c12899 (.ZN (slo__sro_n11829), .A1 (slo__sro_n11830), .A2 (slo__sro_n11831));
AOI21_X4 slo__sro_c12900 (.ZN (slo__sro_n11828), .A (slo__sro_n11829), .B1 (n_6_374), .B2 (n_6_1_940));
NAND2_X1 CLOCK_sgo__sro_c52624 (.ZN (CLOCK_sgo__sro_n48190), .A1 (n_6_1_940), .A2 (n_6_354));
AND2_X1 slo__sro_c12949 (.ZN (slo__sro_n11872), .A1 (CLOCK_opt_ipo_n46137), .A2 (CLOCK_sgo__n46950));
NAND2_X1 CLOCK_slo__sro_c61602 (.ZN (CLOCK_slo__sro_n55930), .A1 (slo__sro_n6239), .A2 (CLOCK_sgo__n46922));
INV_X2 slo__c13065 (.ZN (slo__n11990), .A (n_6_1_361));
INV_X4 opt_ipo_c49464 (.ZN (opt_ipo_n45121), .A (CLOCK_sgo__sro_n47822));
INV_X1 slo__c13083 (.ZN (slo__n12005), .A (n_6_1_1089));
INV_X2 slo__c13095 (.ZN (slo__n12014), .A (slo__sro_n9138));
AND2_X1 slo__sro_c12975 (.ZN (slo__sro_n11889), .A1 (n_6_2352), .A2 (n_6_1_448));
INV_X1 CLOCK_slo__c52927 (.ZN (slo__sro_n15108), .A (CLOCK_slo__n48430));
INV_X1 slo__c13174 (.ZN (slo__n12071), .A (n_6_1_697));
NAND2_X1 slo__sro_c13222 (.ZN (slo__sro_n12111), .A1 (slo__sro_n12112), .A2 (slo__sro_n12113));
BUF_X32 slo__c13007 (.Z (slo__n11938), .A (Multiplier[6]));
AOI21_X2 slo__sro_c13223 (.ZN (slo__sro_n12110), .A (slo__sro_n12111), .B1 (n_6_581), .B2 (n_6_1_799));
NAND2_X1 slo__sro_c13346 (.ZN (slo__sro_n12227), .A1 (CLOCK_opt_ipo_n45978), .A2 (n_6_1_343));
NAND2_X1 slo__sro_c13347 (.ZN (slo__sro_n12226), .A1 (n_6_1415), .A2 (slo___n23229));
INV_X2 slo__L1_c1_c32893 (.ZN (slo__sro_n8179), .A (slo__n29395));
INV_X2 slo__c13309 (.ZN (slo__n12190), .A (slo__sro_n19436));
NAND2_X1 slo__sro_c13348 (.ZN (slo__sro_n12225), .A1 (slo__sro_n12226), .A2 (slo__sro_n12227));
AOI21_X2 slo__sro_c13349 (.ZN (slo__sro_n12224), .A (slo__sro_n12225), .B1 (n_6_1447), .B2 (n_6_1_345));
NAND2_X1 slo__sro_c38246 (.ZN (slo__sro_n34608), .A1 (n_6_410), .A2 (n_6_1_904));
INV_X1 slo__sro_c13378 (.ZN (slo__sro_n12256), .A (slo__sro_n12257));
AOI221_X2 slo__sro_c13379 (.ZN (slo__sro_n12255), .A (slo__sro_n12256), .B1 (n_6_741)
    , .B2 (n_6_1_730), .C1 (n_6_709), .C2 (n_6_1_729));
AOI221_X2 slo__sro_c13580 (.ZN (n_6_1_960), .A (slo__sro_n12409), .B1 (n_6_275), .B2 (n_6_1_974)
    , .C1 (n_6_307), .C2 (n_6_1_975));
NAND2_X1 slo__sro_c13688 (.ZN (slo__sro_n12492), .A1 (n_6_922), .A2 (slo___n23367));
NAND2_X1 slo__sro_c13689 (.ZN (slo__sro_n12491), .A1 (slo__sro_n12492), .A2 (slo__sro_n12493));
AOI21_X2 slo__sro_c13690 (.ZN (slo__sro_n12490), .A (slo__sro_n12491), .B1 (n_6_954), .B2 (n_6_1_625));
INV_X1 slo__sro_c13704 (.ZN (slo__sro_n12507), .A (n_6_1_658));
NOR2_X1 slo__sro_c13705 (.ZN (slo__sro_n12506), .A1 (slo__sro_n12508), .A2 (slo__sro_n12507));
INV_X1 CLOCK_slo__sro_c55025 (.ZN (CLOCK_slo__sro_n50321), .A (slo__sro_n8966));
NAND2_X1 slo__sro_c13725 (.ZN (slo__sro_n12525), .A1 (n_6_2663), .A2 (n_6_1_798));
INV_X1 slo__sro_c13726 (.ZN (slo__sro_n12524), .A (slo__sro_n12525));
AOI221_X1 slo__sro_c13727 (.ZN (n_6_1_794), .A (slo__sro_n12524), .B1 (n_6_604), .B2 (n_6_1_799)
    , .C1 (n_6_636), .C2 (n_6_1_800));
NAND2_X1 slo__sro_c13763 (.ZN (slo__sro_n12556), .A1 (slo__sro_n12557), .A2 (slo__sro_n12558));
AOI21_X2 slo__sro_c13764 (.ZN (n_6_1_829), .A (slo__sro_n12556), .B1 (n_6_572), .B2 (n_6_1_835));
NAND2_X1 slo__sro_c13778 (.ZN (slo__sro_n12570), .A1 (n_6_1304), .A2 (n_6_1_414));
NAND2_X1 slo__sro_c13779 (.ZN (slo__sro_n12569), .A1 (slo__sro_n12570), .A2 (slo__sro_n12571));
AOI21_X2 slo__sro_c13780 (.ZN (slo__sro_n12568), .A (slo__sro_n12569), .B1 (n_6_1336), .B2 (slo___n43257));
AOI222_X2 slo__sro_c14126 (.ZN (slo__sro_n12865), .A1 (n_6_593), .A2 (n_6_1_799), .B1 (n_6_625)
    , .B2 (n_6_1_800), .C1 (n_6_2652), .C2 (n_6_1_798));
NAND2_X1 slo__sro_c13983 (.ZN (slo__sro_n12746), .A1 (n_6_2216), .A2 (n_6_1_308));
INV_X2 slo__c13821 (.ZN (slo__n12606), .A (n_6_1_649));
NAND2_X1 slo__sro_c13984 (.ZN (slo__sro_n12745), .A1 (n_6_1487), .A2 (n_6_1_309));
NAND2_X1 slo__sro_c13985 (.ZN (slo__sro_n12744), .A1 (slo__sro_n12745), .A2 (slo__sro_n12746));
AOI21_X2 slo__sro_c13986 (.ZN (slo__sro_n12743), .A (slo__sro_n12744), .B1 (n_6_1519), .B2 (slo___n23247));
INV_X2 slo__c14064 (.ZN (slo__n12818), .A (n_6_1_824));
INV_X1 slo__c14101 (.ZN (slo__n12843), .A (n_6_1_325));
INV_X1 slo___L1_c1_c14398 (.ZN (slo___n13099), .A (CLOCK_slo__xsl_n57029));
AOI222_X2 slo__sro_c14154 (.ZN (n_6_1_713), .A1 (n_6_721), .A2 (n_6_1_729), .B1 (n_6_753)
    , .B2 (n_6_1_730), .C1 (n_6_2590), .C2 (n_6_1_728));
NAND2_X1 slo__sro_c14192 (.ZN (slo__sro_n12925), .A1 (n_6_1550), .A2 (n_6_1_274));
NAND2_X1 slo__sro_c14193 (.ZN (slo__sro_n12924), .A1 (slo__sro_n12925), .A2 (slo__sro_n12926));
NAND2_X1 CLOCK_slo__sro_c66519 (.ZN (CLOCK_slo__sro_n59962), .A1 (n_6_304), .A2 (n_6_1_975));
INV_X1 opt_ipo_c27187 (.ZN (opt_ipo_n23804), .A (slo__sro_n32716));
CLKBUF_X1 slo__c14345 (.Z (slo__n13053), .A (n_6_2011));
AND2_X1 slo__sro_c14236 (.ZN (slo__sro_n12963), .A1 (n_6_2656), .A2 (n_6_1_798));
AOI21_X1 slo__sro_c25230 (.ZN (slo__sro_n22026), .A (slo__sro_n9390), .B1 (n_6_1603), .B2 (slo___n23215));
INV_X1 slo__c14256 (.ZN (slo__n12976), .A (slo__sro_n19970));
NAND2_X1 CLOCK_slo__sro_c66072 (.ZN (CLOCK_slo__sro_n59551), .A1 (n_6_1_343), .A2 (n_6_2233));
NAND2_X1 slo__sro_c15142 (.ZN (slo__sro_n13701), .A1 (slo__sro_n13702), .A2 (slo__sro_n13703));
NAND2_X1 slo__sro_c14557 (.ZN (slo__sro_n13235), .A1 (n_6_2135), .A2 (n_6_1_203));
BUF_X32 drc_ipo_c29984 (.Z (drc_ipo_n26610), .A (Multiplier[15]));
INV_X2 slo__c14460 (.ZN (slo__n13153), .A (CLOCK_sgo__sro_n47592));
NAND2_X1 slo__sro_c14679 (.ZN (slo__sro_n13335), .A1 (n_6_2222), .A2 (n_6_1_308));
NAND2_X1 slo__sro_c14558 (.ZN (slo__sro_n13234), .A1 (n_6_1691), .A2 (n_6_1_204));
NAND2_X1 slo__sro_c14559 (.ZN (slo__sro_n13233), .A1 (slo__sro_n13234), .A2 (slo__sro_n13235));
AOI21_X2 slo__sro_c14560 (.ZN (slo__sro_n13232), .A (slo__sro_n13233), .B1 (n_6_1723), .B2 (slo___n23407));
NAND2_X1 slo__sro_c14680 (.ZN (slo__sro_n13334), .A1 (n_6_1493), .A2 (n_6_1_309));
INV_X1 slo__c14643 (.ZN (slo__n13303), .A (slo__sro_n31234));
NAND2_X1 slo__sro_c14681 (.ZN (slo__sro_n13333), .A1 (slo__sro_n13334), .A2 (slo__sro_n13335));
AND2_X1 slo__sro_c14661 (.ZN (slo__sro_n13318), .A1 (n_6_2162), .A2 (n_6_1_238));
NAND2_X1 slo__sro_c25552 (.ZN (slo__sro_n22328), .A1 (n_6_2897), .A2 (slo__n13799));
NAND2_X2 slo__sro_c14706 (.ZN (slo__sro_n13355), .A1 (slo__sro_n13356), .A2 (slo__sro_n13357));
AOI21_X4 slo__sro_c14707 (.ZN (slo__sro_n13354), .A (slo__sro_n13355), .B1 (n_6_1783), .B2 (CLOCK_sgo__n48020));
NAND2_X2 slo__sro_c14721 (.ZN (slo__sro_n13371), .A1 (n_6_1788), .A2 (CLOCK_sgo__n48020));
NAND2_X4 slo__sro_c14722 (.ZN (slo__sro_n13370), .A1 (slo__sro_n13371), .A2 (slo__sro_n13372));
AND2_X1 CLOCK_slo__sro_c63591 (.ZN (CLOCK_slo__sro_n57490), .A1 (n_6_81), .A2 (n_6_1_1079));
NAND2_X1 slo__sro_c14737 (.ZN (slo__sro_n13384), .A1 (n_6_1710), .A2 (slo___n23407));
NAND2_X2 slo__sro_c14738 (.ZN (slo__sro_n13383), .A1 (slo__sro_n13384), .A2 (slo__sro_n13385));
AOI21_X4 slo__sro_c14739 (.ZN (slo__sro_n13382), .A (slo__sro_n13383), .B1 (n_6_1678), .B2 (slo___n23239));
INV_X2 slo__c14751 (.ZN (slo__n13394), .A (slo__n15804));
NAND2_X1 slo__sro_c14841 (.ZN (slo__sro_n13473), .A1 (n_6_1360), .A2 (n_6_1_379));
NAND2_X1 slo__sro_c14842 (.ZN (slo__sro_n13472), .A1 (slo__sro_n13473), .A2 (slo__sro_n13474));
INV_X1 slo__c14780 (.ZN (slo__n13417), .A (slo__sro_n21662));
NAND2_X1 CLOCK_slo__sro_c53530 (.ZN (CLOCK_slo__sro_n48978), .A1 (n_6_2057), .A2 (n_6_1_133));
AND2_X1 slo__sro_c14907 (.ZN (slo__sro_n13522), .A1 (n_6_2747), .A2 (CLOCK_sgo__n46934));
INV_X1 slo__c14804 (.ZN (slo__n13438), .A (n_6_1_811));
NAND2_X1 slo__sro_c41271 (.ZN (slo__sro_n37388), .A1 (slo__sro_n37389), .A2 (slo__sro_n37390));
INV_X1 slo__c14920 (.ZN (slo__n13528), .A (CLOCK_slo__sro_n49772));
AOI21_X4 CLOCK_slo__sro_c53837 (.ZN (n_6_1_511), .A (CLOCK_slo__sro_n49242), .B1 (n_6_1145), .B2 (slo___n23268));
NAND2_X1 slo__sro_c15140 (.ZN (slo__sro_n13703), .A1 (n_6_2360), .A2 (n_6_1_483));
INV_X1 slo__c15040 (.ZN (slo__n13621), .A (n_6_1_646));
NAND2_X1 slo__sro_c15141 (.ZN (slo__sro_n13702), .A1 (n_6_1156), .A2 (slo___n23364));
AOI21_X2 slo__sro_c15143 (.ZN (slo__sro_n13700), .A (slo__sro_n13701), .B1 (n_6_1188), .B2 (slo___n23466));
INV_X1 slo__c14971 (.ZN (slo__n13570), .A (n_6_1_488));
INV_X2 slo__c15026 (.ZN (slo__n13610), .A (n_6_1_684));
INV_X1 slo__c14882 (.ZN (slo__n13501), .A (slo__sro_n36476));
INV_X1 slo__c19939 (.ZN (slo__n17556), .A (n_6_1_676));
NAND2_X1 slo__sro_c15182 (.ZN (slo__sro_n13738), .A1 (slo__sro_n17353), .A2 (slo__sro_n13740));
NAND2_X1 CLOCK_slo__sro_c57683 (.ZN (CLOCK_slo__sro_n52593), .A1 (CLOCK_slo__sro_n52594), .A2 (CLOCK_slo__sro_n52595));
INV_X2 slo__c15171 (.ZN (slo__n13728), .A (slo__sro_n6817));
INV_X2 slo__L1_c1_c32954 (.ZN (n_6_1_757), .A (slo__n29454));
AND2_X1 CLOCK_slo__sro_c65942 (.ZN (CLOCK_slo__sro_n59437), .A1 (n_6_2256), .A2 (n_6_1_343));
INV_X1 slo__c15328 (.ZN (slo__n13851), .A (slo__sro_n6519));
INV_X2 slo__c15309 (.ZN (slo__n13838), .A (slo__sro_n37482));
INV_X1 slo__c15402 (.ZN (slo__n13910), .A (n_6_1_777));
INV_X1 slo__c15262 (.ZN (n_6_1_1074), .A (slo__sro_n37221));
AOI21_X1 CLOCK_slo__sro_c68984 (.ZN (CLOCK_slo__sro_n62128), .A (CLOCK_slo__sro_n62129)
    , .B1 (n_6_205), .B2 (n_6_1_1009));
BUF_X32 drc_ipo_c29956 (.Z (drc_ipo_n26579), .A (n_6_20));
NAND2_X1 slo__sro_c15458 (.ZN (slo__sro_n13954), .A1 (n_6_621), .A2 (n_6_1_800));
BUF_X4 drc_ipo_c29969 (.Z (drc_ipo_n26592), .A (n_6_10));
INV_X1 slo__c15347 (.ZN (slo__n13864), .A (slo__sro_n39888));
INV_X1 slo__c15392 (.ZN (slo__n13903), .A (slo__sro_n6229));
NAND2_X1 slo__sro_c15459 (.ZN (slo__sro_n13953), .A1 (slo__sro_n13954), .A2 (slo__sro_n13955));
AOI21_X2 slo__sro_c15460 (.ZN (n_6_1_779), .A (slo__sro_n13953), .B1 (n_6_589), .B2 (n_6_1_799));
NAND2_X1 CLOCK_sgo__sro_c51983 (.ZN (CLOCK_sgo__sro_n47664), .A1 (slo___n23215), .A2 (n_6_1608));
INV_X2 slo__c15550 (.ZN (slo__n14026), .A (n_6_1_632));
INV_X1 slo__c15540 (.ZN (slo__n14019), .A (slo__sro_n7037));
INV_X1 slo__c15564 (.ZN (slo__n14037), .A (slo__sro_n20259));
INV_X2 slo__c15434 (.ZN (slo__n13933), .A (slo__sro_n21560));
NAND2_X1 slo__sro_c15618 (.ZN (slo__sro_n14083), .A1 (n_6_1428), .A2 (slo___n23229));
NAND2_X1 slo__sro_c15619 (.ZN (slo__sro_n14082), .A1 (slo__sro_n14083), .A2 (slo__sro_n14084));
AOI222_X2 slo__sro_c15520 (.ZN (n_6_1_998), .A1 (n_6_246), .A2 (n_6_1_1010), .B1 (n_6_214)
    , .B2 (n_6_1_1009), .C1 (n_6_2843), .C2 (CLOCK_sgo__n46950));
INV_X1 slo__c15634 (.ZN (slo__n14095), .A (slo__sro_n6191));
NAND2_X1 slo__sro_c15725 (.ZN (slo__sro_n14165), .A1 (n_6_1686), .A2 (n_6_1_204));
INV_X1 slo__c15646 (.ZN (slo__n14104), .A (n_6_1_120));
INV_X1 slo__c15658 (.ZN (slo__n14113), .A (n_6_1_627));
INV_X2 slo__c15674 (.ZN (slo__n14126), .A (n_6_1_630));
NAND2_X1 slo__sro_c15726 (.ZN (slo__sro_n14164), .A1 (slo__sro_n14165), .A2 (slo__sro_n14166));
AOI21_X1 slo__sro_c15727 (.ZN (slo__sro_n14163), .A (slo__sro_n14164), .B1 (n_6_1718), .B2 (slo___n23407));
NAND2_X2 slo__sro_c39308 (.ZN (slo__sro_n35616), .A1 (slo__sro_n35617), .A2 (slo__sro_n35618));
INV_X1 slo__c15697 (.ZN (slo__n14143), .A (n_6_1_233));
INV_X2 slo__c15774 (.ZN (slo__n14207), .A (n_6_1_259));
NAND2_X1 CLOCK_sgo__sro_c51345 (.ZN (CLOCK_sgo__sro_n47136), .A1 (slo___n13086), .A2 (n_6_1_378));
INV_X1 slo__sro_c15855 (.ZN (slo__sro_n14274), .A (slo__sro_n14275));
AOI221_X1 slo__sro_c15856 (.ZN (n_6_1_1035), .A (slo__sro_n14274), .B1 (n_6_184), .B2 (n_6_1_1045)
    , .C1 (n_6_152), .C2 (n_6_1_1044));
AOI21_X2 slo__c15910 (.ZN (slo__n14340), .A (slo__sro_n9008), .B1 (n_6_67), .B2 (n_6_1_1079));
AOI222_X2 slo__sro_c16140 (.ZN (n_6_1_712), .A1 (n_6_720), .A2 (n_6_1_729), .B1 (n_6_752)
    , .B2 (n_6_1_730), .C1 (n_6_2589), .C2 (n_6_1_728));
INV_X2 slo__c16058 (.ZN (slo__n14465), .A (slo__sro_n4784));
INV_X1 slo__sro_c32502 (.ZN (slo__sro_n29018), .A (slo__sro_n29019));
AND2_X1 CLOCK_slo__sro_c70258 (.ZN (n_6_1_956), .A1 (CLOCK_slo__sro_n63268), .A2 (CLOCK_slo__sro_n63269));
INV_X2 slo__c16088 (.ZN (slo__n14486), .A (n_6_1_756));
NAND2_X1 slo__sro_c16125 (.ZN (slo__sro_n14524), .A1 (n_6_358), .A2 (n_6_1_940));
NAND2_X2 slo__sro_c16126 (.ZN (slo__sro_n14523), .A1 (slo__sro_n14524), .A2 (slo__sro_n14525));
AOI21_X4 slo__sro_c16127 (.ZN (slo__sro_n14522), .A (slo__sro_n14523), .B1 (n_6_326), .B2 (n_6_1_939));
AOI222_X2 slo__sro_c16299 (.ZN (n_6_1_124), .A1 (n_6_1847), .A2 (n_6_1_135), .B1 (n_6_1815)
    , .B2 (n_6_1_134), .C1 (n_6_2069), .C2 (n_6_1_133));
INV_X1 slo__c16264 (.ZN (slo__n14633), .A (n_6_1_1034));
INV_X1 slo__c16274 (.ZN (slo__n14640), .A (n_6_1_324));
INV_X2 slo__c16284 (.ZN (slo__n14647), .A (slo__sro_n19751));
INV_X1 slo__c16328 (.ZN (slo__n14684), .A (CLOCK_slo__sro_n48812));
INV_X1 slo__c16254 (.ZN (slo__n14626), .A (slo__sro_n21314));
INV_X1 slo__c16338 (.ZN (slo__n14691), .A (slo__sro_n21676));
NAND2_X1 slo__sro_c30535 (.ZN (slo__sro_n27160), .A1 (n_6_2041), .A2 (n_6_1_98));
INV_X2 slo__c43674 (.ZN (slo__n39406), .A (n_6_1_330));
AOI222_X2 slo__sro_c16407 (.ZN (slo__sro_n14742), .A1 (n_6_1744), .A2 (n_6_1_169)
    , .B1 (n_6_1776), .B2 (CLOCK_sgo__n48020), .C1 (n_6_2093), .C2 (n_6_1_168));
INV_X1 slo__c16442 (.ZN (slo__n14771), .A (n_6_1_155));
INV_X2 slo__c16434 (.ZN (slo__n14766), .A (slo__sro_n13278));
INV_X1 slo__c16365 (.ZN (slo__n14709), .A (n_6_1_711));
NAND2_X1 slo__sro_c16537 (.ZN (slo__sro_n14855), .A1 (slo__sro_n14856), .A2 (slo__sro_n14857));
INV_X2 slo__c41061 (.ZN (slo__n37202), .A (slo__sro_n27860));
INV_X1 slo__c16586 (.ZN (slo__n14899), .A (CLOCK_slo__sro_n54647));
INV_X2 slo__c16578 (.ZN (slo__n14894), .A (n_6_1_968));
NAND2_X1 CLOCK_slo__sro_c69771 (.ZN (CLOCK_slo__sro_n62841), .A1 (CLOCK_slo__sro_n62842), .A2 (CLOCK_slo__sro_n62843));
INV_X2 slo__c16635 (.ZN (slo__n14942), .A (slo__sro_n34034));
BUF_X32 drc_ipo_c29968 (.Z (drc_ipo_n26591), .A (n_6_9));
INV_X1 slo__c16645 (.ZN (slo__n14949), .A (slo__n39180));
AOI222_X2 slo__sro_c16742 (.ZN (slo__sro_n15043), .A1 (n_6_547), .A2 (n_6_1_835), .B1 (n_6_515)
    , .B2 (n_6_1_834), .C1 (slo__sro_n15108), .C2 (CLOCK_sgo__n46922));
CLKBUF_X1 spw__L1_c1_c76597 (.Z (n_6_2856), .A (spw__n68416));
NAND2_X2 slo__sro_c16665 (.ZN (CLOCK_slo__n60839), .A1 (CLOCK_opt_ipo_n45730), .A2 (hfn_ipo_n35));
INV_X1 slo__sro_c16814 (.ZN (slo__sro_n15109), .A (slo__sro_n15110));
AOI221_X1 slo__sro_c16815 (.ZN (CLOCK_slo__n48430), .A (slo__sro_n15109), .B1 (n_6_484)
    , .B2 (n_6_1_870), .C1 (n_6_452), .C2 (n_6_1_869));
NAND2_X1 slo__sro_c16897 (.ZN (slo__sro_n15185), .A1 (n_6_2191), .A2 (n_6_1_273));
INV_X1 slo__c16873 (.ZN (slo__n15162), .A (n_6_1_967));
NAND2_X1 slo__sro_c16898 (.ZN (slo__sro_n15184), .A1 (n_6_1557), .A2 (n_6_1_274));
INV_X1 slo__sro_c16850 (.ZN (slo__sro_n15145), .A (n_6_2767));
INV_X1 slo__sro_c16851 (.ZN (slo__sro_n15144), .A (CLOCK_sgo__n46937));
NOR2_X1 slo__sro_c16852 (.ZN (slo__sro_n15143), .A1 (slo__sro_n15145), .A2 (slo__sro_n15144));
INV_X1 slo__sro_c25889 (.ZN (slo__sro_n22625), .A (n_6_2846));
INV_X2 CLOCK_slo__c55530 (.ZN (n_6_1_995), .A (CLOCK_slo__n50780));
NAND2_X1 CLOCK_slo__sro_c56661 (.ZN (CLOCK_slo__sro_n51766), .A1 (n_6_829), .A2 (n_6_1_695));
INV_X1 slo__c16989 (.ZN (slo__n15246), .A (slo__sro_n27391));
AND2_X1 slo__sro_c17109 (.ZN (slo__sro_n15343), .A1 (n_6_2158), .A2 (n_6_1_238));
INV_X2 slo__L1_c1_c39510 (.ZN (slo__n35802), .A (slo__sro_n37819));
NAND2_X1 slo__sro_c17154 (.ZN (slo__sro_n15382), .A1 (n_6_2773), .A2 (CLOCK_sgo__n46937));
INV_X1 slo__c17029 (.ZN (slo__n15271), .A (n_6_1_919));
NAND2_X1 slo__sro_c17155 (.ZN (slo__sro_n15381), .A1 (n_6_366), .A2 (n_6_1_940));
NAND2_X1 slo__sro_c17156 (.ZN (slo__sro_n15380), .A1 (slo__sro_n15381), .A2 (slo__sro_n15382));
AOI21_X1 slo__sro_c17157 (.ZN (n_6_1_920), .A (slo__sro_n15380), .B1 (n_6_334), .B2 (n_6_1_939));
INV_X1 slo__c17210 (.ZN (slo__n15420), .A (n_6_1_223));
INV_X2 slo__c17243 (.ZN (slo__n15443), .A (slo__sro_n27138));
INV_X1 slo__c16981 (.ZN (slo__n15241), .A (n_6_1_923));
NAND2_X1 slo__sro_c17277 (.ZN (slo__sro_n15471), .A1 (n_6_1665), .A2 (n_6_1_204));
NAND2_X1 slo__sro_c17278 (.ZN (slo__sro_n15470), .A1 (slo__sro_n15472), .A2 (slo__sro_n15471));
AOI21_X2 slo__sro_c17279 (.ZN (n_6_1_172), .A (slo__sro_n15470), .B1 (n_6_1697), .B2 (slo___n23407));
NAND2_X1 slo__sro_c17293 (.ZN (slo__sro_n15484), .A1 (n_6_1610), .A2 (slo___n23215));
NAND2_X1 slo__sro_c17294 (.ZN (slo__sro_n15483), .A1 (slo__sro_n15484), .A2 (slo__sro_n15485));
AOI21_X1 slo__sro_c17295 (.ZN (slo__sro_n15482), .A (slo__sro_n15483), .B1 (n_6_1642), .B2 (drc_ipo_n26601));
AOI221_X2 slo__sro_c17399 (.ZN (slo__sro_n15586), .A (slo__sro_n15587), .B1 (n_6_278)
    , .B2 (n_6_1_974), .C1 (n_6_310), .C2 (n_6_1_975));
AOI222_X1 slo__sro_c17353 (.ZN (slo__n28071), .A1 (n_6_1839), .A2 (n_6_1_135), .B1 (n_6_1807)
    , .B2 (slo___n43254), .C1 (n_6_2061), .C2 (n_6_1_133));
NAND2_X4 slo__sro_c17499 (.ZN (slo__sro_n15670), .A1 (n_6_1560), .A2 (n_6_1_274));
BUF_X32 slo__c30082 (.Z (slo__n26713), .A (drc_ipo_n26595));
AOI21_X4 slo__sro_c17501 (.ZN (slo__sro_n15668), .A (slo__sro_n15669), .B1 (n_6_1592), .B2 (slo___n23244));
INV_X2 CLOCK_slo__mro_c57198 (.ZN (CLOCK_slo__mro_n52174), .A (n_6_934));
INV_X1 CLOCK_slo__mro_c57199 (.ZN (slo__sro_n42343), .A (n_6_1_625));
AOI21_X2 slo__sro_c17517 (.ZN (slo__sro_n15684), .A (slo__sro_n15685), .B1 (n_6_1591), .B2 (slo___n23244));
NAND2_X1 slo__sro_c17531 (.ZN (slo__sro_n15702), .A1 (n_6_1545), .A2 (n_6_1_274));
NAND2_X1 slo__sro_c17532 (.ZN (slo__sro_n15701), .A1 (slo__sro_n15702), .A2 (slo__sro_n15703));
AOI21_X1 slo__sro_c17533 (.ZN (slo__sro_n15700), .A (slo__sro_n15701), .B1 (n_6_1577), .B2 (slo___n23244));
AND2_X1 slo__sro_c17629 (.ZN (slo__sro_n15779), .A1 (n_6_2257), .A2 (n_6_1_343));
NAND2_X1 slo__sro_c24646 (.ZN (slo__sro_n21500), .A1 (n_6_2896), .A2 (slo__n13799));
AND2_X1 slo__sro_c17647 (.ZN (slo__sro_n15796), .A1 (n_6_2117), .A2 (n_6_1_203));
AOI222_X1 CLOCK_slo__sro_c63123 (.ZN (n_6_1_993), .A1 (n_6_241), .A2 (n_6_1_1010)
    , .B1 (n_6_209), .B2 (n_6_1_1009), .C1 (slo___n8281), .C2 (CLOCK_sgo__n46950));
NAND2_X1 slo__sro_c17691 (.ZN (slo__sro_n15832), .A1 (opt_ipo_n24707), .A2 (n_6_1_168));
INV_X1 slo__c17682 (.ZN (slo__n15821), .A (n_6_1_143));
NAND2_X1 slo__sro_c17693 (.ZN (slo__sro_n15830), .A1 (slo__sro_n15831), .A2 (slo__sro_n15832));
AOI21_X2 slo__sro_c17694 (.ZN (CLOCK_slo__n48906), .A (slo__sro_n15830), .B1 (n_6_1774), .B2 (CLOCK_sgo__n48020));
INV_X2 slo__c17587 (.ZN (slo__n15745), .A (slo__sro_n14742));
AOI21_X1 slo__sro_c17857 (.ZN (slo__sro_n15955), .A (n_6_1_132), .B1 (n_6_1821), .B2 (n_6_1_134));
INV_X2 slo__c17792 (.ZN (slo__n15903), .A (slo__sro_n27726));
INV_X1 slo__c17756 (.ZN (slo__n15879), .A (n_6_1_121));
AND2_X2 slo__sro_c17858 (.ZN (n_6_1_130), .A1 (slo__sro_n15956), .A2 (slo__sro_n15955));
INV_X2 slo__c17936 (.ZN (slo__n16022), .A (n_6_1_160));
INV_X1 slo__c17744 (.ZN (slo__n15870), .A (n_6_1_162));
INV_X2 slo__c17887 (.ZN (slo__n15976), .A (n_6_1_909));
INV_X1 slo__c17777 (.ZN (slo__n15894), .A (n_6_1_268));
INV_X1 slo__c17877 (.ZN (slo__n15969), .A (slo__sro_n10769));
INV_X2 slo__c17998 (.ZN (slo__n16063), .A (n_6_1_127));
NAND2_X1 slo__sro_c17911 (.ZN (slo__sro_n16003), .A1 (n_6_1_168), .A2 (n_6_2098));
NAND2_X1 slo__sro_c17912 (.ZN (slo__sro_n16002), .A1 (n_6_1749), .A2 (n_6_1_169));
NAND2_X1 slo__sro_c17913 (.ZN (slo__sro_n16001), .A1 (slo__sro_n16002), .A2 (slo__sro_n16003));
INV_X1 slo__c17831 (.ZN (slo__n15930), .A (n_6_1_267));
INV_X1 CLOCK_slo__sro_c56308 (.ZN (CLOCK_slo__sro_n51475), .A (n_6_1_202));
NAND2_X1 slo__sro_c18164 (.ZN (slo__sro_n16183), .A1 (n_6_2647), .A2 (n_6_1_798));
AOI21_X2 CLOCK_slo__sro_c63142 (.ZN (n_6_1_809), .A (CLOCK_slo__sro_n57154), .B1 (n_6_520), .B2 (n_6_1_834));
NAND2_X1 slo__sro_c18165 (.ZN (slo__sro_n16182), .A1 (n_6_620), .A2 (n_6_1_800));
NAND2_X1 slo__sro_c18166 (.ZN (slo__sro_n16181), .A1 (slo__sro_n16182), .A2 (slo__sro_n16183));
INV_X1 slo__c18130 (.ZN (slo__n16152), .A (slo__sro_n5794));
AOI21_X1 slo__sro_c18167 (.ZN (slo__sro_n16180), .A (slo__sro_n16181), .B1 (n_6_588), .B2 (n_6_1_799));
NAND2_X1 slo__sro_c18207 (.ZN (slo__sro_n16216), .A1 (slo__sro_n16217), .A2 (slo__sro_n16218));
NAND2_X1 slo__sro_c33404 (.ZN (slo__sro_n29880), .A1 (slo__sro_n4752), .A2 (slo__sro_n29881));
AOI21_X1 slo__sro_c18208 (.ZN (slo__sro_n16215), .A (slo__sro_n16216), .B1 (n_6_136), .B2 (n_6_1_1044));
NAND2_X1 CLOCK_sgo__sro_c51501 (.ZN (CLOCK_sgo__sro_n47262), .A1 (n_6_1_274), .A2 (n_6_1554));
NOR2_X1 slo__sro_c35288 (.ZN (slo__sro_n31655), .A1 (slo__sro_n31657), .A2 (slo__sro_n31656));
NAND2_X1 slo__sro_c35794 (.ZN (slo__sro_n32140), .A1 (opt_ipo_n24326), .A2 (CLOCK_sgo__n46937));
INV_X1 slo__c18274 (.ZN (slo__n16267), .A (n_6_1_511));
INV_X2 slo__c18293 (.ZN (slo__n16280), .A (n_6_1_825));
INV_X1 slo__c18524 (.ZN (slo__n16450), .A (n_6_1_396));
INV_X2 slo__c18389 (.ZN (slo__n16348), .A (slo__sro_n6038));
BUF_X8 drc_ipo_c29972 (.Z (drc_ipo_n26595), .A (slo__n3834));
INV_X1 slo__c18451 (.ZN (slo__n16392), .A (n_6_1_828));
AOI222_X2 slo__sro_c19075 (.ZN (slo__sro_n16886), .A1 (n_6_1195), .A2 (slo___n23466)
    , .B1 (n_6_1163), .B2 (slo___n23364), .C1 (n_6_2367), .C2 (n_6_1_483));
INV_X1 slo__c18955 (.ZN (slo__n16796), .A (n_6_1_827));
INV_X1 slo__c18381 (.ZN (slo__n16343), .A (n_6_1_717));
INV_X1 slo__c18622 (.ZN (slo__n16524), .A (slo__sro_n4615));
BUF_X32 slo__c18721 (.Z (slo__n16608), .A (slo__n38599));
INV_X1 slo__c18630 (.ZN (slo__n16529), .A (slo__sro_n9701));
INV_X4 slo__c18663 (.ZN (slo__n16550), .A (sgo__sro_n1599));
INV_X1 slo__c18481 (.ZN (slo__n16413), .A (slo__sro_n11215));
INV_X2 slo__c18673 (.ZN (slo__n16557), .A (n_6_1_894));
INV_X1 slo__c19272 (.ZN (slo__n17041), .A (n_6_1_513));
INV_X1 slo__c18897 (.ZN (slo__n16747), .A (n_6_1_359));
AOI221_X2 slo__sro_c30283 (.ZN (slo__sro_n11578), .A (slo__sro_n26911), .B1 (n_6_215)
    , .B2 (n_6_1_1009), .C1 (n_6_247), .C2 (n_6_1_1010));
BUF_X32 slo__c18694 (.Z (slo__n16572), .A (CLOCK_slo___n64878));
INV_X2 slo__c18850 (.ZN (slo__n16706), .A (CLOCK_slo__sro_n55687));
INV_X2 slo__c18947 (.ZN (slo__n16791), .A (sgo__sro_n1557));
INV_X1 slo__sro_c19290 (.ZN (slo__sro_n17058), .A (n_6_2845));
INV_X2 slo__c18927 (.ZN (slo__n16774), .A (n_6_1_969));
INV_X1 slo__c19191 (.ZN (slo__n16975), .A (n_6_1_536));
INV_X1 slo__c19060 (.ZN (slo__n16871), .A (slo__sro_n7852));
INV_X1 slo__c19050 (.ZN (slo__n16864), .A (CLOCK_slo__sro_n53339));
AOI21_X2 slo__sro_c19105 (.ZN (slo__sro_n16910), .A (slo__sro_n5225), .B1 (n_6_1252), .B2 (slo___n23274));
INV_X1 slo__sro_c19291 (.ZN (slo__sro_n17057), .A (CLOCK_sgo__n46950));
INV_X1 slo__c19245 (.ZN (slo__n17020), .A (slo__sro_n9559));
NOR2_X1 slo__sro_c19292 (.ZN (slo__sro_n17056), .A1 (slo__sro_n17058), .A2 (slo__sro_n17057));
AOI221_X2 slo__sro_c19293 (.ZN (n_6_1_1000), .A (slo__sro_n17056), .B1 (n_6_248), .B2 (n_6_1_1010)
    , .C1 (n_6_216), .C2 (n_6_1_1009));
NAND2_X1 slo__sro_c19312 (.ZN (slo__sro_n17076), .A1 (n_6_2546), .A2 (n_6_1_693));
INV_X1 slo__sro_c19313 (.ZN (slo__sro_n17075), .A (slo__sro_n17076));
AOI221_X1 slo__sro_c19314 (.ZN (slo__sro_n17074), .A (slo__sro_n17075), .B1 (n_6_804)
    , .B2 (n_6_1_695), .C1 (n_6_772), .C2 (n_6_1_694));
INV_X1 slo__sro_c19546 (.ZN (slo__sro_n17256), .A (n_6_2859));
INV_X1 slo__c19506 (.ZN (slo__n17214), .A (n_6_1_549));
INV_X1 slo__sro_c19547 (.ZN (slo__sro_n17255), .A (CLOCK_sgo__n46945));
NAND2_X1 slo__sro_c19532 (.ZN (slo__sro_n17239), .A1 (slo__sro_n17240), .A2 (slo__sro_n17241));
NOR2_X1 slo__sro_c19548 (.ZN (slo__sro_n17254), .A1 (slo__sro_n17256), .A2 (slo__sro_n17255));
NAND2_X1 slo__sro_c19530 (.ZN (slo__sro_n17241), .A1 (n_6_2898), .A2 (slo__n13799));
NAND2_X1 slo__sro_c19531 (.ZN (slo__sro_n17240), .A1 (n_6_1_1080), .A2 (n_6_111));
AOI21_X1 slo__sro_c19533 (.ZN (slo__sro_n17238), .A (slo__sro_n17239), .B1 (n_6_79), .B2 (n_6_1_1079));
NAND2_X1 slo__sro_c34643 (.ZN (slo__sro_n31051), .A1 (slo__sro_n31052), .A2 (slo__sro_n31053));
AOI221_X1 CLOCK_slo__sro_c66623 (.ZN (slo__sro_n39513), .A (CLOCK_slo__sro_n60053)
    , .B1 (n_6_1766), .B2 (n_6_1_170), .C1 (n_6_1734), .C2 (n_6_1_169));
INV_X1 slo__c19592 (.ZN (slo__n17290), .A (CLOCK_slo__sro_n56057));
AOI222_X2 slo__sro_c19644 (.ZN (slo__sro_n17330), .A1 (n_6_1205), .A2 (slo___n23466)
    , .B1 (n_6_1173), .B2 (slo___n23364), .C1 (n_6_2377), .C2 (n_6_1_483));
INV_X1 slo__c19785 (.ZN (slo__n17435), .A (n_6_1_475));
INV_X1 slo__c19710 (.ZN (slo__n17378), .A (n_6_1_369));
AND2_X1 slo__sro_c19992 (.ZN (slo__sro_n17598), .A1 (n_6_2413), .A2 (n_6_1_518));
CLKBUF_X1 spw__L1_c1_c76463 (.Z (n_6_1993), .A (spw__n68268));
AOI221_X2 CLOCK_slo__sro_c65722 (.ZN (slo__sro_n9845), .A (CLOCK_slo__sro_n59232)
    , .B1 (n_6_1097), .B2 (slo___n23277), .C1 (n_6_1129), .C2 (slo___n23268));
NAND2_X4 slo__sro_c20055 (.ZN (slo__sro_n17647), .A1 (slo__sro_n17648), .A2 (slo__sro_n17649));
INV_X2 slo__c19961 (.ZN (slo__n17575), .A (n_6_1_575));
INV_X1 slo__c19737 (.ZN (slo__n17399), .A (slo__sro_n7435));
NAND2_X1 slo__sro_c20053 (.ZN (slo__sro_n17649), .A1 (n_6_1_483), .A2 (n_6_2381));
INV_X2 slo__c19763 (.ZN (slo__n17416), .A (n_6_1_371));
NAND2_X2 slo__sro_c20054 (.ZN (slo__sro_n17648), .A1 (n_6_1177), .A2 (slo___n23364));
INV_X2 slo__c20017 (.ZN (slo__n17619), .A (slo__n17737));
AOI21_X2 slo__sro_c20056 (.ZN (slo__sro_n17646), .A (slo__sro_n17647), .B1 (n_6_1209), .B2 (slo___n23466));
AND2_X2 slo__sro_c20231 (.ZN (n_6_1_707), .A1 (slo__sro_n17781), .A2 (slo__sro_n17782));
INV_X1 slo__c20087 (.ZN (slo__n17671), .A (n_6_1_158));
AND2_X1 slo__sro_c20190 (.ZN (slo__sro_n17753), .A1 (n_6_2415), .A2 (n_6_1_518));
INV_X1 slo__c20099 (.ZN (slo__n17680), .A (n_6_1_123));
NAND2_X1 CLOCK_slo__sro_c53694 (.ZN (CLOCK_slo__sro_n49121), .A1 (n_6_2490), .A2 (n_6_1_623));
AOI222_X1 slo__sro_c40655 (.ZN (spw__n66802), .A1 (n_6_775), .A2 (n_6_1_694), .B1 (n_6_807)
    , .B2 (n_6_1_695), .C1 (n_6_2549), .C2 (n_6_1_693));
INV_X2 slo__c20181 (.ZN (slo__n17744), .A (slo__sro_n32044));
AOI221_X2 slo__sro_c20203 (.ZN (n_6_1_548), .A (slo__sro_n17761), .B1 (n_6_1051), .B2 (n_6_1_554)
    , .C1 (n_6_1083), .C2 (slo___n23457));
NAND2_X1 slo__sro_c20229 (.ZN (slo__sro_n17782), .A1 (n_6_715), .A2 (n_6_1_729));
AOI21_X1 slo__sro_c20230 (.ZN (slo__sro_n17781), .A (slo__sro_n5332), .B1 (n_6_747), .B2 (n_6_1_730));
NOR2_X1 slo__sro_c45434 (.ZN (slo__sro_n40960), .A1 (slo__sro_n40962), .A2 (slo__sro_n40961));
INV_X1 slo__c20282 (.ZN (slo__n17821), .A (slo__sro_n19997));
AOI221_X2 CLOCK_slo__sro_c56362 (.ZN (CLOCK_slo__sro_n51511), .A (CLOCK_slo__sro_n51512)
    , .B1 (n_6_919), .B2 (slo___n23367), .C1 (n_6_951), .C2 (n_6_1_625));
INV_X1 slo__c20422 (.ZN (slo__n17921), .A (slo__sro_n13262));
NAND2_X1 CLOCK_slo__sro_c56402 (.ZN (CLOCK_slo__sro_n51543), .A1 (n_6_908), .A2 (slo___n23367));
AOI21_X4 slo__sro_c20464 (.ZN (n_6_1_562), .A (slo__sro_n17951), .B1 (n_6_966), .B2 (slo___n23232));
NAND2_X1 slo__sro_c21047 (.ZN (slo__sro_n18406), .A1 (n_6_1_238), .A2 (n_6_2153));
INV_X2 slo__c20545 (.ZN (slo__n18019), .A (CLOCK_sgo__sro_n47798));
INV_X1 slo__c20452 (.ZN (slo__n17942), .A (n_6_1_1004));
NAND2_X1 slo__sro_c20571 (.ZN (slo__sro_n18044), .A1 (slo___n16361), .A2 (n_6_1_448));
AOI221_X2 slo__sro_c20573 (.ZN (slo__sro_n18042), .A (slo__sro_n18043), .B1 (n_6_1249)
    , .B2 (slo___n23274), .C1 (n_6_1217), .C2 (slo___n23359));
INV_X2 slo__c20623 (.ZN (slo__n18079), .A (slo__sro_n7583));
CLKBUF_X1 spw__L1_c1_c77590 (.Z (spw__n69100), .A (spw__n69101));
INV_X1 slo__c20894 (.ZN (slo__n18286), .A (n_6_1_563));
INV_X1 slo__c20911 (.ZN (slo__n18297), .A (n_6_1_949));
NAND2_X1 slo__sro_c20725 (.ZN (slo__sro_n18156), .A1 (n_6_2174), .A2 (n_6_1_273));
INV_X2 slo__c20681 (.ZN (slo__n18122), .A (n_6_1_187));
NAND2_X1 slo__sro_c20726 (.ZN (slo__sro_n18155), .A1 (n_6_1540), .A2 (n_6_1_274));
NAND2_X1 slo__sro_c20727 (.ZN (slo__sro_n18154), .A1 (slo__sro_n18155), .A2 (slo__sro_n18156));
NAND2_X2 CLOCK_slo__sro_c56799 (.ZN (CLOCK_slo__sro_n51887), .A1 (n_6_1511), .A2 (slo___n23247));
INV_X2 slo__c20759 (.ZN (slo__n18178), .A (n_6_1_457));
AOI21_X2 CLOCK_slo__sro_c63885 (.ZN (CLOCK_slo__sro_n57699), .A (CLOCK_slo__sro_n57700)
    , .B1 (n_6_1598), .B2 (slo___n23244));
NAND2_X1 CLOCK_slo__sro_c57758 (.ZN (CLOCK_slo__sro_n52671), .A1 (n_6_1_588), .A2 (n_6_2471));
INV_X1 slo__c20954 (.ZN (slo__n18328), .A (slo__sro_n22132));
NAND2_X1 slo__sro_c21049 (.ZN (slo__sro_n18404), .A1 (slo__sro_n18405), .A2 (slo__sro_n18406));
AOI21_X1 slo__sro_c21050 (.ZN (slo__sro_n18403), .A (slo__sro_n18404), .B1 (n_6_1646), .B2 (drc_ipo_n26601));
INV_X1 slo__c21127 (.ZN (slo__n18465), .A (n_6_1_950));
INV_X1 slo__sro_c21143 (.ZN (slo__sro_n18480), .A (slo__sro_n18481));
AOI221_X2 slo__sro_c21144 (.ZN (n_6_1_879), .A (slo__sro_n18480), .B1 (n_6_424), .B2 (n_6_1_905)
    , .C1 (n_6_392), .C2 (n_6_1_904));
AND2_X1 CLOCK_slo__sro_c53217 (.ZN (CLOCK_slo__sro_n48699), .A1 (n_6_1700), .A2 (slo___n23407));
AND2_X1 slo__sro_c21780 (.ZN (slo__sro_n18951), .A1 (n_6_2144), .A2 (n_6_1_238));
BUF_X4 drc_ipo_c29965 (.Z (drc_ipo_n26588), .A (n_6_12));
INV_X1 slo__c21195 (.ZN (slo__n18523), .A (CLOCK_slo__sro_n51132));
INV_X2 slo__c21459 (.ZN (slo__n18727), .A (n_6_1_1072));
INV_X1 slo__c21467 (.ZN (slo__n18732), .A (n_6_1_1037));
INV_X1 slo__c21325 (.ZN (slo__n18626), .A (n_6_1_1038));
INV_X1 slo__c21361 (.ZN (slo__n18653), .A (slo__sro_n40769));
INV_X1 slo__c21521 (.ZN (slo__n18771), .A (n_6_1_915));
INV_X1 slo__c21513 (.ZN (slo__n18766), .A (slo__sro_n29674));
INV_X1 slo__c21529 (.ZN (slo__n18776), .A (n_6_1_951));
AND2_X1 slo__sro_c21652 (.ZN (slo__sro_n18863), .A1 (n_6_2815), .A2 (n_6_1_973));
INV_X1 slo__sro_c35286 (.ZN (slo__sro_n31657), .A (n_6_2855));
INV_X1 CLOCK_slo__sro_c56489 (.ZN (CLOCK_slo__sro_n51621), .A (slo__sro_n36933));
INV_X1 slo__c21771 (.ZN (slo__n18942), .A (n_6_1_706));
INV_X2 slo__c21673 (.ZN (slo__n18877), .A (slo__sro_n11828));
INV_X1 slo__c21637 (.ZN (slo__n18848), .A (slo__sro_n6790));
NAND2_X1 slo__sro_c21939 (.ZN (slo__sro_n19079), .A1 (slo___n19182), .A2 (n_6_1_798));
INV_X1 slo__c21930 (.ZN (slo__n19067), .A (slo__sro_n17693));
INV_X1 slo__c21812 (.ZN (slo__n18973), .A (n_6_1_703));
INV_X1 slo__c21839 (.ZN (slo__n18991), .A (slo__sro_n4312));
INV_X4 slo__c21827 (.ZN (slo__n18982), .A (slo__sro_n13354));
NAND2_X1 slo__sro_c21940 (.ZN (slo__sro_n19078), .A1 (n_6_1_799), .A2 (n_6_595));
NAND2_X1 slo__sro_c21941 (.ZN (slo__sro_n19077), .A1 (slo__sro_n19078), .A2 (slo__sro_n19079));
NAND2_X1 slo__sro_c21872 (.ZN (slo__sro_n19027), .A1 (n_6_2178), .A2 (n_6_1_273));
NAND2_X1 slo__sro_c21873 (.ZN (slo__sro_n19026), .A1 (n_6_1544), .A2 (n_6_1_274));
NAND2_X1 slo__sro_c21874 (.ZN (slo__sro_n19025), .A1 (slo__sro_n19026), .A2 (slo__sro_n19027));
AOI21_X1 slo__sro_c21875 (.ZN (slo__sro_n19024), .A (slo__sro_n19025), .B1 (n_6_1576), .B2 (slo___n23244));
INV_X1 CLOCK_sgo__L1_c1_c51291 (.ZN (CLOCK_sgo__n47093), .A (CLOCK_sgo__n47094));
BUF_X4 drc_ipo_c29971 (.Z (drc_ipo_n26594), .A (n_6_6));
INV_X1 slo__c21971 (.ZN (slo__n19102), .A (n_6_1_819));
AOI21_X2 slo__sro_c22326 (.ZN (n_6_1_711), .A (slo__sro_n19349), .B1 (n_6_751), .B2 (n_6_1_730));
INV_X1 slo__c22229 (.ZN (slo__n19282), .A (CLOCK_slo__sro_n60275));
NAND2_X1 slo__sro_c22363 (.ZN (slo__sro_n19384), .A1 (n_6_282), .A2 (n_6_1_974));
NAND2_X1 slo__sro_c22324 (.ZN (slo__sro_n19350), .A1 (n_6_1_729), .A2 (n_6_719));
INV_X2 slo__c22081 (.ZN (slo__n19179), .A (n_6_1_496));
NAND2_X1 slo__sro_c22325 (.ZN (slo__sro_n19349), .A1 (slo__sro_n19350), .A2 (slo__sro_n19351));
INV_X1 slo__c22187 (.ZN (slo__n19255), .A (n_6_1_712));
INV_X1 slo__c22282 (.ZN (slo__n19320), .A (slo__sro_n3748));
NAND2_X1 slo__sro_c22364 (.ZN (slo__sro_n19383), .A1 (slo__sro_n19384), .A2 (slo__sro_n19385));
AOI21_X2 slo__sro_c22365 (.ZN (n_6_1_967), .A (slo__sro_n19383), .B1 (n_6_314), .B2 (n_6_1_975));
NAND2_X1 slo__sro_c22404 (.ZN (slo__sro_n19422), .A1 (n_6_1300), .A2 (n_6_1_414));
NAND2_X1 slo__sro_c22405 (.ZN (slo__sro_n19421), .A1 (slo__sro_n19422), .A2 (slo__sro_n19423));
AOI21_X4 slo__sro_c22406 (.ZN (slo__sro_n19420), .A (slo__sro_n19421), .B1 (n_6_1332), .B2 (slo___n43257));
NAND2_X1 slo__sro_c22420 (.ZN (slo__sro_n19438), .A1 (n_6_1_764), .A2 (n_6_647));
NAND2_X2 slo__sro_c22421 (.ZN (slo__sro_n19437), .A1 (slo__sro_n19438), .A2 (slo__sro_n19439));
AOI21_X2 slo__sro_c22422 (.ZN (slo__sro_n19436), .A (slo__sro_n19437), .B1 (n_6_679), .B2 (n_6_1_765));
AND2_X1 slo__sro_c46788 (.ZN (slo__sro_n42332), .A1 (slo___n13777), .A2 (n_6_1_728));
NAND2_X1 slo__sro_c22539 (.ZN (slo__sro_n19546), .A1 (n_6_1_448), .A2 (opt_ipo_n23778));
NAND2_X1 CLOCK_slo__sro_c56403 (.ZN (CLOCK_slo__sro_n51542), .A1 (CLOCK_slo__sro_n51543), .A2 (CLOCK_slo__sro_n51544));
AOI21_X1 CLOCK_slo__sro_c56404 (.ZN (CLOCK_slo__sro_n51541), .A (CLOCK_slo__sro_n51542)
    , .B1 (n_6_940), .B2 (n_6_1_625));
AOI21_X2 slo__sro_c22542 (.ZN (slo__sro_n19543), .A (slo__sro_n19544), .B1 (n_6_1222), .B2 (slo___n23359));
NAND2_X1 slo__sro_c22565 (.ZN (slo__sro_n19568), .A1 (slo__sro_n19569), .A2 (slo__sro_n19570));
AOI21_X2 slo__sro_c22566 (.ZN (slo__sro_n19567), .A (slo__sro_n19568), .B1 (n_6_1338), .B2 (slo___n43257));
NAND2_X1 slo__sro_c22758 (.ZN (slo__sro_n19753), .A1 (n_6_1435), .A2 (slo___n23229));
NAND2_X1 slo__sro_c22759 (.ZN (slo__sro_n19752), .A1 (slo__sro_n19753), .A2 (slo__sro_n19754));
INV_X1 slo__sro_c22997 (.ZN (slo__sro_n19972), .A (n_6_1_588));
AND2_X1 slo__sro_c22625 (.ZN (slo__sro_n19628), .A1 (n_6_2225), .A2 (n_6_1_308));
NAND2_X1 CLOCK_sgo__sro_c51534 (.ZN (CLOCK_sgo__sro_n47286), .A1 (CLOCK_sgo__sro_n47287), .A2 (slo__sro_n28564));
AND2_X1 slo__sro_c22731 (.ZN (slo__sro_n19728), .A1 (n_6_2501), .A2 (n_6_1_623));
AND2_X1 CLOCK_slo__sro_c70042 (.ZN (CLOCK_slo__sro_n63090), .A1 (n_6_493), .A2 (n_6_1_870));
AND2_X1 slo__sro_c22849 (.ZN (slo__sro_n19839), .A1 (n_6_2875), .A2 (CLOCK_sgo__n46945));
NAND2_X1 slo__sro_c22757 (.ZN (slo__sro_n19754), .A1 (n_6_2259), .A2 (n_6_1_343));
NAND2_X1 slo__sro_c22814 (.ZN (slo__sro_n19806), .A1 (slo__sro_n19807), .A2 (slo__sro_n19808));
AOI21_X2 slo__sro_c22815 (.ZN (slo__sro_n19805), .A (slo__sro_n19806), .B1 (n_6_529), .B2 (n_6_1_834));
AOI221_X2 slo__sro_c22850 (.ZN (n_6_1_1034), .A (slo__sro_n19839), .B1 (n_6_183), .B2 (n_6_1_1045)
    , .C1 (n_6_151), .C2 (n_6_1_1044));
NAND2_X1 slo__sro_c22671 (.ZN (slo__sro_n19676), .A1 (n_6_2253), .A2 (n_6_1_343));
NAND2_X2 slo__sro_c22672 (.ZN (slo__sro_n19675), .A1 (n_6_1429), .A2 (slo___n23229));
NAND2_X2 slo__sro_c22673 (.ZN (slo__sro_n19674), .A1 (slo__sro_n19675), .A2 (slo__sro_n19676));
AOI21_X2 slo__sro_c22674 (.ZN (slo__sro_n19673), .A (slo__sro_n19674), .B1 (n_6_1461), .B2 (n_6_1_345));
AOI221_X2 slo__sro_c22999 (.ZN (slo__sro_n19970), .A (slo__sro_n19971), .B1 (n_6_972)
    , .B2 (slo___n23232), .C1 (n_6_1004), .C2 (slo___n23218));
NAND2_X1 slo__sro_c22984 (.ZN (slo__sro_n19960), .A1 (n_6_2462), .A2 (n_6_1_588));
INV_X1 slo__sro_c22985 (.ZN (slo__sro_n19959), .A (slo__sro_n19960));
AOI221_X2 slo__sro_c22986 (.ZN (slo__sro_n19958), .A (slo__sro_n19959), .B1 (n_6_973)
    , .B2 (slo___n23232), .C1 (n_6_1005), .C2 (slo___n23218));
NAND2_X1 slo__sro_c22914 (.ZN (slo__sro_n19897), .A1 (n_6_2716), .A2 (n_6_1_868));
NAND2_X1 slo__sro_c22915 (.ZN (slo__sro_n19896), .A1 (n_6_467), .A2 (n_6_1_869));
NAND2_X1 slo__sro_c22916 (.ZN (slo__sro_n19895), .A1 (slo__sro_n19896), .A2 (slo__sro_n19897));
AOI21_X2 slo__sro_c22917 (.ZN (slo__sro_n19894), .A (slo__sro_n19895), .B1 (n_6_499), .B2 (n_6_1_870));
INV_X2 CLOCK_slo__c55736 (.ZN (n_6_1_782), .A (CLOCK_slo__n50956));
NAND2_X1 slo__sro_c23102 (.ZN (slo__sro_n20067), .A1 (n_6_1_939), .A2 (n_6_343));
NAND2_X1 slo__sro_c23103 (.ZN (slo__sro_n20066), .A1 (slo__sro_n20067), .A2 (slo__sro_n20068));
AOI21_X2 slo__sro_c23104 (.ZN (n_6_1_929), .A (slo__sro_n20066), .B1 (n_6_375), .B2 (n_6_1_940));
AOI222_X2 slo__sro_c43619 (.ZN (slo__sro_n39363), .A1 (n_6_1865), .A2 (CLOCK_sgo__n48011)
    , .B1 (n_6_1897), .B2 (n_6_1_100), .C1 (n_6_2024), .C2 (n_6_1_98));
NAND2_X1 slo__sro_c23087 (.ZN (slo__sro_n20058), .A1 (n_6_2770), .A2 (CLOCK_sgo__n46937));
NAND2_X1 slo__sro_c23088 (.ZN (slo__sro_n20057), .A1 (n_6_1_940), .A2 (n_6_363));
NAND2_X1 slo__sro_c23089 (.ZN (slo__sro_n20056), .A1 (slo__sro_n20057), .A2 (slo__sro_n20058));
AOI21_X1 slo__sro_c23090 (.ZN (n_6_1_917), .A (slo__sro_n20056), .B1 (n_6_331), .B2 (n_6_1_939));
NAND2_X2 CLOCK_sgo__sro_c52162 (.ZN (CLOCK_sgo__sro_n47800), .A1 (n_6_1371), .A2 (n_6_1_379));
NAND2_X1 slo__sro_c23315 (.ZN (slo__sro_n20260), .A1 (slo__sro_n20261), .A2 (slo__sro_n20262));
AOI21_X1 slo__sro_c23316 (.ZN (slo__sro_n20259), .A (slo__sro_n20260), .B1 (n_6_944), .B2 (n_6_1_625));
NAND2_X1 CLOCK_slo__sro_c56940 (.ZN (CLOCK_slo__sro_n51980), .A1 (CLOCK_slo__sro_n51981), .A2 (CLOCK_slo__sro_n51982));
NAND2_X1 slo__sro_c23341 (.ZN (slo__sro_n20288), .A1 (n_6_2334), .A2 (n_6_1_448));
AND2_X1 slo__sro_c23172 (.ZN (slo__sro_n20127), .A1 (n_6_2204), .A2 (n_6_1_308));
AND2_X1 slo__sro_c36160 (.ZN (slo__sro_n32485), .A1 (n_6_853), .A2 (slo___n23463));
NAND2_X1 slo__sro_c23343 (.ZN (slo__sro_n20286), .A1 (slo__sro_n20287), .A2 (slo__sro_n20288));
AOI21_X1 slo__sro_c23344 (.ZN (slo__sro_n20285), .A (slo__sro_n20286), .B1 (n_6_1225), .B2 (slo___n23359));
AOI21_X2 slo__sro_c23381 (.ZN (slo__sro_n20321), .A (slo__sro_n20322), .B1 (n_6_1132), .B2 (slo___n23268));
INV_X1 slo__sro_c23457 (.ZN (slo__sro_n20395), .A (n_6_1_378));
NOR2_X1 slo__sro_c23458 (.ZN (slo__sro_n20394), .A1 (slo__sro_n20396), .A2 (slo__sro_n20395));
NAND2_X1 CLOCK_slo__sro_c53508 (.ZN (CLOCK_slo__sro_n48960), .A1 (n_6_2212), .A2 (n_6_1_308));
BUF_X2 slo__c34167 (.Z (slo__n30589), .A (sgo__n711));
INV_X1 slo__mro_c36917 (.ZN (slo__mro_n33269), .A (hfn_ipo_n35));
NAND2_X1 slo__mro_c36918 (.ZN (slo__mro_n33268), .A1 (n_6_1981), .A2 (n_6_1_65));
NAND2_X1 slo__sro_c23545 (.ZN (slo__sro_n20475), .A1 (n_6_2203), .A2 (n_6_1_308));
NAND2_X1 slo__sro_c23546 (.ZN (slo__sro_n20474), .A1 (n_6_1474), .A2 (n_6_1_309));
NAND2_X1 slo__sro_c23547 (.ZN (slo__sro_n20473), .A1 (slo__sro_n20474), .A2 (slo__sro_n20475));
AOI21_X2 slo__sro_c23548 (.ZN (slo__sro_n20472), .A (slo__sro_n20473), .B1 (n_6_1506), .B2 (slo___n23247));
NAND2_X1 slo__sro_c23640 (.ZN (slo__sro_n20568), .A1 (n_6_2486), .A2 (n_6_1_623));
NAND2_X1 CLOCK_sgo__sro_c51364 (.ZN (CLOCK_sgo__sro_n47149), .A1 (n_6_739), .A2 (n_6_1_730));
BUF_X1 slo___L1_c47634 (.Z (slo___n43254), .A (n_6_1_134));
NOR2_X1 slo__sro_c23688 (.ZN (slo__sro_n20613), .A1 (slo__sro_n20615), .A2 (slo__sro_n20614));
AOI221_X2 slo__sro_c23689 (.ZN (slo__sro_n20612), .A (slo__sro_n20613), .B1 (n_6_250)
    , .B2 (n_6_1_1010), .C1 (n_6_218), .C2 (n_6_1_1009));
NAND2_X1 slo__sro_c35858 (.ZN (slo__sro_n32204), .A1 (n_6_1_168), .A2 (n_6_2103));
NAND2_X1 slo__sro_c23760 (.ZN (slo__sro_n20682), .A1 (n_6_1303), .A2 (n_6_1_414));
NAND2_X2 slo__sro_c23761 (.ZN (slo__sro_n20681), .A1 (slo__sro_n20682), .A2 (slo__sro_n20683));
AOI21_X4 slo__sro_c23762 (.ZN (slo__sro_n20680), .A (slo__sro_n20681), .B1 (n_6_1335), .B2 (slo___n43257));
NAND2_X1 slo__sro_c23822 (.ZN (slo__sro_n20735), .A1 (n_6_2164), .A2 (n_6_1_238));
INV_X1 slo__sro_c23823 (.ZN (slo__sro_n20734), .A (slo__sro_n20735));
AOI221_X2 slo__sro_c23824 (.ZN (n_6_1_231), .A (slo__sro_n20734), .B1 (n_6_1625), .B2 (slo___n23215)
    , .C1 (n_6_1657), .C2 (drc_ipo_n26601));
NOR2_X1 slo__sro_c23915 (.ZN (slo__sro_n20818), .A1 (slo__sro_n20820), .A2 (slo__sro_n20819));
AOI221_X2 slo__sro_c23916 (.ZN (slo__sro_n20817), .A (slo__sro_n20818), .B1 (n_6_594)
    , .B2 (n_6_1_799), .C1 (n_6_626), .C2 (n_6_1_800));
NAND2_X1 slo__sro_c23942 (.ZN (slo__sro_n20847), .A1 (n_6_500), .A2 (n_6_1_870));
NAND2_X1 slo__sro_c23943 (.ZN (slo__sro_n20846), .A1 (n_6_468), .A2 (n_6_1_869));
AND3_X2 slo__sro_c23944 (.ZN (slo__sro_n20845), .A1 (slo__sro_n20846), .A2 (slo__sro_n20848), .A3 (slo__sro_n20847));
NAND2_X1 slo__sro_c23985 (.ZN (slo__sro_n20887), .A1 (slo___n23367), .A2 (n_6_924));
NAND2_X1 slo__sro_c23986 (.ZN (slo__sro_n20886), .A1 (slo__sro_n20887), .A2 (slo__sro_n20888));
AOI21_X2 slo__sro_c23987 (.ZN (slo__sro_n20885), .A (slo__sro_n20886), .B1 (n_6_956), .B2 (n_6_1_625));
INV_X1 slo__sro_c24013 (.ZN (slo__sro_n20915), .A (slo__sro_n5630));
NAND2_X1 slo__sro_c24014 (.ZN (slo__sro_n20914), .A1 (n_6_1238), .A2 (slo___n23359));
NAND2_X1 slo__sro_c24015 (.ZN (slo__sro_n20913), .A1 (slo__sro_n20914), .A2 (slo__sro_n20915));
AOI21_X2 slo__sro_c24016 (.ZN (n_6_1_438), .A (slo__sro_n20913), .B1 (n_6_1270), .B2 (slo___n23274));
AND2_X1 CLOCK_slo__sro_c63353 (.ZN (CLOCK_slo__sro_n57315), .A1 (n_6_1756), .A2 (slo___n23430));
NAND2_X1 slo__sro_c24125 (.ZN (slo__sro_n21012), .A1 (n_6_633), .A2 (n_6_1_800));
AOI21_X1 slo__sro_c24126 (.ZN (slo__sro_n21011), .A (slo__sro_n4176), .B1 (n_6_601), .B2 (n_6_1_799));
AND2_X1 slo__sro_c24127 (.ZN (n_6_1_791), .A1 (slo__sro_n21011), .A2 (slo__sro_n21012));
NAND2_X2 slo__sro_c24453 (.ZN (slo__sro_n21316), .A1 (n_6_1_905), .A2 (n_6_440));
NAND2_X2 slo__sro_c24454 (.ZN (slo__sro_n21315), .A1 (slo__sro_n21316), .A2 (slo__sro_n21317));
AOI21_X2 slo__sro_c24455 (.ZN (slo__sro_n21314), .A (slo__sro_n21315), .B1 (n_6_408), .B2 (n_6_1_904));
NAND2_X1 slo__sro_c24082 (.ZN (slo__sro_n20974), .A1 (CLOCK_sgo__n46945), .A2 (n_6_2865));
AND2_X1 CLOCK_slo__sro_c69753 (.ZN (CLOCK_slo__sro_n62823), .A1 (CLOCK_slo__sro_n62825), .A2 (CLOCK_slo__sro_n62824));
NAND2_X1 CLOCK_slo__sro_c55601 (.ZN (CLOCK_slo__sro_n50841), .A1 (n_6_302), .A2 (n_6_1_975));
NAND2_X1 slo__sro_c24486 (.ZN (slo__sro_n21348), .A1 (n_6_849), .A2 (slo___n23463));
NAND2_X1 slo__sro_c24487 (.ZN (slo__sro_n21347), .A1 (slo__sro_n21348), .A2 (slo__sro_n21349));
AOI21_X1 slo__sro_c24488 (.ZN (slo__sro_n21346), .A (slo__sro_n21347), .B1 (n_6_881), .B2 (n_6_1_660));
NAND2_X1 slo__sro_c24521 (.ZN (slo__sro_n21382), .A1 (n_6_1_273), .A2 (n_6_2189));
NAND2_X1 slo__sro_c24522 (.ZN (slo__sro_n21381), .A1 (n_6_1_274), .A2 (n_6_1555));
NAND2_X1 slo__sro_c24523 (.ZN (slo__sro_n21380), .A1 (slo__sro_n21381), .A2 (slo__sro_n21382));
AOI21_X2 slo__sro_c24524 (.ZN (n_6_1_260), .A (slo__sro_n21380), .B1 (n_6_1587), .B2 (slo___n23244));
AOI21_X4 slo__sro_c24584 (.ZN (slo__sro_n21436), .A (slo__sro_n21437), .B1 (n_6_1465), .B2 (n_6_1_345));
NAND2_X1 slo__sro_c24647 (.ZN (slo__sro_n21499), .A1 (n_6_109), .A2 (n_6_1_1080));
NAND2_X1 slo__sro_c24648 (.ZN (slo__sro_n21498), .A1 (slo__sro_n21499), .A2 (slo__sro_n21500));
AOI21_X1 slo__sro_c24649 (.ZN (n_6_1_1059), .A (slo__sro_n21498), .B1 (n_6_77), .B2 (n_6_1_1079));
NAND2_X1 CLOCK_slo__sro_c55077 (.ZN (CLOCK_slo__sro_n50364), .A1 (n_6_1_693), .A2 (n_6_2556));
NAND2_X1 slo__sro_c24792 (.ZN (slo__sro_n21634), .A1 (n_6_786), .A2 (n_6_1_694));
AND2_X1 slo__sro_c24761 (.ZN (slo__sro_n21603), .A1 (n_6_2313), .A2 (n_6_1_413));
INV_X1 slo__sro_c45409 (.ZN (slo__sro_n40939), .A (n_6_2336));
AND3_X1 slo__sro_c24794 (.ZN (slo__sro_n21632), .A1 (slo__sro_n21633), .A2 (slo__sro_n21635), .A3 (slo__sro_n21634));
NAND2_X1 slo__sro_c24828 (.ZN (slo__sro_n21664), .A1 (n_6_933), .A2 (n_6_1_625));
NAND2_X1 slo__sro_c24829 (.ZN (slo__sro_n21663), .A1 (slo__sro_n21664), .A2 (slo__sro_n21665));
AOI21_X2 slo__sro_c24830 (.ZN (slo__sro_n21662), .A (slo__sro_n21663), .B1 (n_6_901), .B2 (slo___n23367));
NAND2_X1 CLOCK_slo__sro_c71927 (.ZN (CLOCK_slo__sro_n64638), .A1 (n_6_1896), .A2 (n_6_1_100));
AOI21_X2 CLOCK_sgo__sro_c51751 (.ZN (n_6_1_163), .A (CLOCK_sgo__sro_n47468), .B1 (n_6_1787), .B2 (CLOCK_sgo__n48020));
BUF_X4 drc_ipo_c29963 (.Z (drc_ipo_n26586), .A (n_6_14));
NAND2_X1 slo__sro_c24927 (.ZN (slo__sro_n21755), .A1 (n_6_1_940), .A2 (n_6_359));
NAND2_X1 slo__sro_c24928 (.ZN (slo__sro_n21754), .A1 (slo__sro_n21755), .A2 (slo__sro_n8245));
AOI21_X2 slo__sro_c24929 (.ZN (slo__sro_n21753), .A (slo__sro_n21754), .B1 (n_6_327), .B2 (n_6_1_939));
NAND2_X1 CLOCK_slo__sro_c65839 (.ZN (CLOCK_slo__sro_n59344), .A1 (n_6_946), .A2 (n_6_1_625));
NAND2_X1 slo__sro_c24975 (.ZN (slo__sro_n21797), .A1 (n_6_2642), .A2 (n_6_1_798));
NAND2_X1 slo__sro_c24976 (.ZN (slo__sro_n21796), .A1 (n_6_615), .A2 (n_6_1_800));
NAND2_X1 slo__sro_c24977 (.ZN (slo__sro_n21795), .A1 (slo__sro_n21796), .A2 (slo__sro_n21797));
AOI21_X2 slo__sro_c24978 (.ZN (n_6_1_773), .A (slo__sro_n21795), .B1 (n_6_583), .B2 (n_6_1_799));
AND2_X1 slo__sro_c25144 (.ZN (slo__sro_n21940), .A1 (slo__sro_n21941), .A2 (slo__sro_n21942));
INV_X1 slo__sro_c25231 (.ZN (slo__sro_n22025), .A (slo__sro_n22026));
AOI21_X2 slo__sro_c25232 (.ZN (slo__sro_n22024), .A (slo__sro_n22025), .B1 (n_6_1635), .B2 (drc_ipo_n26601));
NAND2_X2 slo__sro_c25321 (.ZN (slo__sro_n22112), .A1 (n_6_1_764), .A2 (n_6_662));
NAND2_X1 slo__sro_c25322 (.ZN (slo__sro_n22111), .A1 (slo__sro_n22112), .A2 (slo__sro_n22113));
AOI21_X2 slo__sro_c25323 (.ZN (slo__sro_n22110), .A (slo__sro_n22111), .B1 (n_6_694), .B2 (n_6_1_765));
INV_X2 slo__sro_c25343 (.ZN (slo__sro_n22133), .A (slo__sro_n22134));
AOI21_X4 slo__sro_c25344 (.ZN (slo__sro_n22132), .A (slo__sro_n22133), .B1 (n_6_1655), .B2 (drc_ipo_n26601));
NAND2_X1 slo__sro_c25553 (.ZN (slo__sro_n22327), .A1 (n_6_1_1080), .A2 (n_6_110));
NAND2_X1 slo__sro_c25554 (.ZN (slo__sro_n22326), .A1 (slo__sro_n22327), .A2 (slo__sro_n22328));
AOI21_X1 slo__sro_c25555 (.ZN (slo__sro_n22325), .A (slo__sro_n22326), .B1 (n_6_78), .B2 (n_6_1_1079));
INV_X1 slo__mro_c36698 (.ZN (slo__mro_n33032), .A (n_6_718));
INV_X1 slo__mro_c36699 (.ZN (slo__mro_n33031), .A (n_6_1_729));
AOI21_X2 slo__sro_c25580 (.ZN (slo__sro_n22347), .A (slo__mro_n33014), .B1 (n_6_328), .B2 (n_6_1_939));
NAND2_X1 slo__sro_c25656 (.ZN (slo__sro_n22417), .A1 (CLOCK_opt_ipo_n45918), .A2 (n_6_1_448));
INV_X1 slo__sro_c25657 (.ZN (slo__sro_n22416), .A (slo__sro_n22417));
AOI221_X2 slo__sro_c25658 (.ZN (slo__sro_n22415), .A (slo__sro_n22416), .B1 (n_6_1248)
    , .B2 (slo___n23274), .C1 (n_6_1216), .C2 (slo___n23359));
INV_X1 slo__sro_c25676 (.ZN (slo__sro_n22432), .A (slo__sro_n22433));
NAND2_X1 CLOCK_slo__sro_c66621 (.ZN (CLOCK_slo__sro_n60054), .A1 (n_6_2083), .A2 (n_6_1_168));
INV_X1 CLOCK_slo__sro_c60611 (.ZN (CLOCK_slo__sro_n55105), .A (n_6_2570));
NAND2_X1 CLOCK_slo__sro_c69410 (.ZN (CLOCK_slo__sro_n62513), .A1 (n_6_1_379), .A2 (n_6_1346));
NAND2_X1 CLOCK_slo__sro_c69411 (.ZN (CLOCK_slo__sro_n62512), .A1 (CLOCK_slo__sro_n62513), .A2 (CLOCK_slo__sro_n58611));
INV_X1 slo__sro_c25809 (.ZN (slo__sro_n22555), .A (slo__sro_n10956));
NAND2_X1 slo__sro_c35697 (.ZN (slo__sro_n32046), .A1 (n_6_931), .A2 (n_6_1_625));
NAND2_X2 slo__sro_c25811 (.ZN (slo__sro_n22553), .A1 (slo__sro_n22554), .A2 (slo__sro_n22555));
AOI21_X2 slo__sro_c25812 (.ZN (n_6_1_930), .A (slo__sro_n22553), .B1 (n_6_376), .B2 (n_6_1_940));
NOR2_X1 slo__sro_c25891 (.ZN (slo__sro_n22623), .A1 (slo__sro_n22625), .A2 (slo__sro_n22624));
NAND2_X1 CLOCK_slo__sro_c58224 (.ZN (CLOCK_slo__sro_n53080), .A1 (slo__n13799), .A2 (n_6_2892));
NAND2_X1 slo__sro_c25952 (.ZN (slo__sro_n22679), .A1 (n_6_2775), .A2 (CLOCK_sgo__n46937));
INV_X1 slo__sro_c25953 (.ZN (slo__sro_n22678), .A (slo__sro_n22679));
AOI221_X1 slo__sro_c25954 (.ZN (slo__sro_n22677), .A (slo__sro_n22678), .B1 (n_6_336)
    , .B2 (n_6_1_939), .C1 (n_6_368), .C2 (n_6_1_940));
AND2_X1 slo__sro_c25978 (.ZN (slo__sro_n22701), .A1 (slo__sro_n22702), .A2 (slo__sro_n22703));
INV_X1 slo__sro_c26011 (.ZN (slo__sro_n22735), .A (slo__sro_n22736));
AOI221_X2 slo__sro_c26012 (.ZN (n_6_1_927), .A (slo__sro_n22735), .B1 (n_6_373), .B2 (n_6_1_940)
    , .C1 (n_6_341), .C2 (n_6_1_939));
NAND2_X1 slo__sro_c26023 (.ZN (slo__sro_n22744), .A1 (n_6_851), .A2 (slo___n23463));
NAND2_X1 slo__sro_c26024 (.ZN (slo__sro_n22743), .A1 (slo__sro_n22744), .A2 (slo__sro_n22745));
AOI21_X2 slo__sro_c26025 (.ZN (n_6_1_645), .A (slo__sro_n22743), .B1 (n_6_883), .B2 (slo___n23451));
INV_X2 slo__sro_c26074 (.ZN (slo__sro_n22781), .A (n_6_280));
NAND2_X1 slo__sro_c26059 (.ZN (slo__sro_n22771), .A1 (CLOCK_slo__n56734), .A2 (CLOCK_sgo__n46937));
NAND2_X1 slo__sro_c26060 (.ZN (slo__sro_n22770), .A1 (n_6_371), .A2 (n_6_1_940));
NAND2_X1 slo__sro_c26061 (.ZN (slo__sro_n22769), .A1 (slo__sro_n22770), .A2 (slo__sro_n22771));
AOI21_X1 slo__sro_c26062 (.ZN (n_6_1_925), .A (slo__sro_n22769), .B1 (n_6_339), .B2 (n_6_1_939));
OAI21_X2 slo__sro_c26076 (.ZN (slo__sro_n22779), .A (slo__sro_n22782), .B1 (slo__sro_n22781), .B2 (slo__sro_n22780));
AOI21_X2 slo__sro_c26077 (.ZN (n_6_1_965), .A (slo__sro_n22779), .B1 (n_6_312), .B2 (n_6_1_975));
INV_X1 slo__sro_c26178 (.ZN (slo__sro_n22874), .A (slo__sro_n22875));
AOI222_X2 slo__sro_c40932 (.ZN (slo__sro_n37092), .A1 (n_6_497), .A2 (n_6_1_870), .B1 (n_6_465)
    , .B2 (n_6_1_869), .C1 (n_6_2714), .C2 (n_6_1_868));
INV_X1 slo__sro_c26281 (.ZN (slo__sro_n22964), .A (slo__sro_n22965));
NAND2_X1 CLOCK_slo__sro_c69831 (.ZN (CLOCK_slo__sro_n62894), .A1 (n_6_156), .A2 (n_6_1_1044));
AND2_X1 slo__sro_c26465 (.ZN (slo__sro_n23125), .A1 (n_6_2240), .A2 (n_6_1_343));
INV_X1 CLOCK_slo__c58782 (.ZN (CLOCK_slo__n53562), .A (slo__sro_n33466));
NAND2_X1 slo__sro_c40763 (.ZN (slo__sro_n36946), .A1 (n_6_2484), .A2 (n_6_1_623));
BUF_X8 slo___L1_c26577 (.Z (slo___n23218), .A (n_6_1_590));
BUF_X1 slo___L1_c26580 (.Z (slo___n23221), .A (CLOCK_sgo__n48011));
BUF_X1 slo___L1_c26585 (.Z (slo___n23226), .A (n_6_1_134));
BUF_X8 slo___L1_c26588 (.Z (slo___n23229), .A (n_6_1_344));
BUF_X8 slo___L1_c26591 (.Z (slo___n23232), .A (n_6_1_589));
BUF_X1 slo___L1_c26594 (.Z (slo___n23235), .A (n_6_1_100));
BUF_X4 drc_ipo_c29950 (.Z (drc_ipo_n26573), .A (n_6_28));
BUF_X1 slo___L1_c26598 (.Z (slo___n23239), .A (n_6_1_204));
BUF_X8 slo___L1_c26603 (.Z (slo___n23244), .A (n_6_1_275));
BUF_X8 slo___L1_c26606 (.Z (slo___n23247), .A (n_6_1_310));
BUF_X8 slo___L1_c26630 (.Z (slo___n23268), .A (n_6_1_520));
BUF_X4 drc_ipo_c29954 (.Z (drc_ipo_n26577), .A (n_6_21));
BUF_X32 slo___L1_c26636 (.Z (slo___n23274), .A (n_6_1_450));
BUF_X8 slo___L1_c26639 (.Z (slo___n23277), .A (n_6_1_519));
BUF_X32 drc_ipo_c29951 (.Z (drc_ipo_n26574), .A (n_6_27));
BUF_X1 slo___L1_c26724 (.Z (slo___n23353), .A (n_6_1_554));
NAND2_X2 CLOCK_slo__mro_c69069 (.ZN (CLOCK_slo__mro_n62208), .A1 (CLOCK_slo__mro_n62209), .A2 (slo__sro_n22580));
INV_X1 slo__c26624 (.ZN (slo__n23263), .A (slo__n23262));
INV_X16 slo__c26625 (.ZN (n_6_1_309), .A (slo__n23263));
BUF_X16 slo___L1_c26730 (.Z (slo___n23359), .A (n_6_1_449));
BUF_X32 slo___L1_c26735 (.Z (slo___n23364), .A (n_6_1_484));
BUF_X32 slo___L1_c26738 (.Z (slo___n23367), .A (n_6_1_624));
BUF_X1 slo___L1_c26778 (.Z (slo___n23404), .A (n_6_1_135));
BUF_X32 slo___L1_c26781 (.Z (slo___n23407), .A (n_6_1_205));
BUF_X1 slo___L1_c26807 (.Z (slo___n23430), .A (n_6_1_169));
BUF_X1 slo___L1_c26831 (.Z (slo___n23451), .A (n_6_1_660));
INV_X1 slo__c26663 (.ZN (slo__n23299), .A (slo__n23298));
INV_X4 slo__c26664 (.ZN (n_6_1_379), .A (slo__n23299));
BUF_X8 drc_ipo_c29952 (.Z (CLOCK_sgo__n47054), .A (n_6_24));
BUF_X8 slo___L1_c26837 (.Z (slo___n23457), .A (n_6_1_555));
NAND2_X1 CLOCK_slo__sro_c68049 (.ZN (CLOCK_slo__sro_n61284), .A1 (slo___n23229), .A2 (n_6_1420));
BUF_X8 slo___L1_c26843 (.Z (slo___n23463), .A (n_6_1_659));
BUF_X32 slo___L1_c26846 (.Z (slo___n23466), .A (n_6_1_485));
BUF_X32 drc_ipo_c29986 (.Z (drc_ipo_n26614), .A (Multiplier[19]));
INV_X1 slo__c26801 (.ZN (slo__n23425), .A (slo__n23424));
INV_X16 slo__c26802 (.ZN (n_6_1_625), .A (slo__n23425));
INV_X1 slo__c26825 (.ZN (slo__n23446), .A (slo__n23445));
INV_X16 slo__c26826 (.ZN (n_6_1_345), .A (slo__n23446));
BUF_X32 drc_ipo_c29987 (.Z (drc_ipo_n26615), .A (Multiplier[20]));
INV_X1 slo__c26772 (.ZN (slo__n23399), .A (slo__n23398));
INV_X16 slo__c26773 (.ZN (n_6_1_380), .A (slo__n23399));
BUF_X32 drc_ipo_c29988 (.Z (drc_ipo_n26616), .A (Multiplier[21]));
BUF_X32 drc_ipo_c29989 (.Z (drc_ipo_n26617), .A (Multiplier[22]));
BUF_X32 drc_ipo_c29990 (.Z (drc_ipo_n26618), .A (Multiplier[23]));
BUF_X32 drc_ipo_c29991 (.Z (drc_ipo_n26620), .A (Multiplier[24]));
BUF_X32 drc_ipo_c29992 (.Z (CLOCK_sgo__n46841), .A (Multiplier[25]));
BUF_X32 drc_ipo_c29993 (.Z (drc_ipo_n26624), .A (Multiplier[28]));
BUF_X32 drc_ipo_c29994 (.Z (drc_ipo_n26625), .A (Multiplier[29]));
NAND2_X1 CLOCK_slo__sro_c69751 (.ZN (CLOCK_slo__sro_n62825), .A1 (n_6_651), .A2 (n_6_1_764));
NAND2_X1 CLOCK_slo__sro_c69770 (.ZN (CLOCK_slo__sro_n62842), .A1 (n_6_298), .A2 (n_6_1_975));
AOI21_X2 CLOCK_slo__sro_c69714 (.ZN (CLOCK_slo__sro_n62783), .A (CLOCK_slo__sro_n62784)
    , .B1 (n_6_878), .B2 (n_6_1_660));
BUF_X2 slo__L19_c20_c30008 (.Z (slo__n26638), .A (slo__n26645));
NAND2_X1 CLOCK_slo__sro_c69713 (.ZN (CLOCK_slo__sro_n62784), .A1 (CLOCK_slo__sro_n62785), .A2 (CLOCK_slo__sro_n62786));
AOI21_X1 CLOCK_slo__sro_c69671 (.ZN (slo__sro_n33562), .A (CLOCK_slo__sro_n62745)
    , .B1 (n_6_491), .B2 (n_6_1_870));
NAND2_X1 CLOCK_slo__sro_c69670 (.ZN (CLOCK_slo__sro_n62745), .A1 (CLOCK_slo__sro_n49069), .A2 (CLOCK_slo__sro_n62746));
NAND2_X1 CLOCK_slo__sro_c69669 (.ZN (CLOCK_slo__sro_n62746), .A1 (n_6_459), .A2 (n_6_1_869));
CLKBUF_X2 spt__c74558 (.Z (n_6_1_47), .A (spt__n66349));
AOI221_X2 CLOCK_slo__sro_c69580 (.ZN (n_6_1_627), .A (CLOCK_slo__sro_n62668), .B1 (n_6_865)
    , .B2 (n_6_1_660), .C1 (n_6_833), .C2 (slo___n23463));
BUF_X1 slo__L12_c13_c30015 (.Z (slo__n26645), .A (slo__n26648));
INV_X1 CLOCK_slo__sro_c69579 (.ZN (CLOCK_slo__sro_n62668), .A (CLOCK_slo__sro_n62669));
NOR2_X2 CLOCK_slo__sro_c69435 (.ZN (CLOCK_slo__sro_n62530), .A1 (CLOCK_slo__sro_n62531), .A2 (slo__sro_n8580));
BUF_X1 slo__L9_c10_c30018 (.Z (slo__n26648), .A (slo__n26654));
NOR2_X4 CLOCK_slo__mro_c69070 (.ZN (slo__sro_n41478), .A1 (CLOCK_slo__mro_n62208), .A2 (slo__sro_n41479));
AND2_X1 CLOCK_slo__sro_c69383 (.ZN (slo__sro_n34126), .A1 (CLOCK_slo__sro_n62489), .A2 (CLOCK_slo__sro_n62488));
NAND2_X1 CLOCK_slo__sro_c68981 (.ZN (CLOCK_slo__sro_n62131), .A1 (CLOCK_sgo__n46950), .A2 (n_6_2834));
AOI21_X1 CLOCK_slo__sro_c68773 (.ZN (n_6_1_90), .A (CLOCK_slo__sro_n61943), .B1 (n_6_1912), .B2 (n_6_1_100));
INV_X2 opt_ipo_c27255 (.ZN (opt_ipo_n23872), .A (sgo__sro_n1213));
NAND2_X1 CLOCK_slo__sro_c68770 (.ZN (CLOCK_slo__sro_n61945), .A1 (n_6_1_98), .A2 (n_6_2039));
AND2_X1 CLOCK_slo__sro_c68174 (.ZN (CLOCK_slo__sro_n61394), .A1 (CLOCK_slo__sro_n61396), .A2 (CLOCK_slo__sro_n61395));
NAND2_X1 CLOCK_slo__sro_c68771 (.ZN (CLOCK_slo__sro_n61944), .A1 (n_6_1880), .A2 (CLOCK_sgo__n48011));
INV_X1 slo__L2_c31_c30028 (.ZN (slo__n26658), .A (n_6_8));
NAND2_X1 CLOCK_slo__sro_c68793 (.ZN (CLOCK_slo__sro_n61962), .A1 (n_6_1200), .A2 (slo___n23466));
BUF_X32 slo__c30174 (.Z (slo__n26805), .A (drc_ipo_n26594));
NAND2_X1 slo__sro_c30633 (.ZN (slo__sro_n27253), .A1 (n_6_2596), .A2 (n_6_1_728));
INV_X1 slo__sro_c30536 (.ZN (slo__sro_n27159), .A (slo__sro_n27160));
NAND2_X1 slo__sro_c30281 (.ZN (slo__sro_n26912), .A1 (n_6_2844), .A2 (CLOCK_sgo__n46950));
AOI21_X4 slo__sro_c30992 (.ZN (slo__sro_n27581), .A (slo__sro_n27582), .B1 (n_6_761), .B2 (n_6_1_730));
NAND2_X1 slo__sro_c30634 (.ZN (slo__sro_n27252), .A1 (n_6_727), .A2 (n_6_1_729));
NAND2_X1 slo__sro_c30635 (.ZN (slo__sro_n27251), .A1 (slo__sro_n27253), .A2 (slo__sro_n27252));
INV_X1 slo__sro_c38245 (.ZN (slo__sro_n34609), .A (slo__sro_n10098));
NAND2_X1 slo__sro_c30755 (.ZN (slo__sro_n27360), .A1 (slo__sro_n27361), .A2 (slo__sro_n27362));
AOI222_X2 CLOCK_slo__sro_c71493 (.ZN (CLOCK_slo__sro_n64272), .A1 (n_6_892), .A2 (slo___n23451)
    , .B1 (n_6_860), .B2 (slo___n23463), .C1 (n_6_2539), .C2 (n_6_1_658));
BUF_X1 slo__L2_c2_c30265 (.Z (slo__n26894), .A (slo__n26895));
INV_X2 slo__L1_c1_c30266 (.ZN (slo__n26895), .A (slo__n26896));
NAND2_X1 slo__sro_c30515 (.ZN (slo__sro_n27140), .A1 (n_6_2097), .A2 (n_6_1_168));
INV_X1 slo__sro_c30753 (.ZN (slo__sro_n27362), .A (slo__sro_n8559));
AOI21_X2 slo__sro_c30636 (.ZN (n_6_1_719), .A (slo__sro_n27251), .B1 (n_6_759), .B2 (n_6_1_730));
AOI21_X2 slo__sro_c30756 (.ZN (slo__sro_n8558), .A (slo__sro_n27360), .B1 (n_6_825), .B2 (n_6_1_695));
AND2_X1 slo__sro_c30789 (.ZN (slo__sro_n27392), .A1 (n_6_2777), .A2 (CLOCK_sgo__n46937));
AOI222_X2 CLOCK_slo__sro_c58520 (.ZN (CLOCK_slo__sro_n53339), .A1 (n_6_311), .A2 (n_6_1_975)
    , .B1 (n_6_279), .B2 (n_6_1_974), .C1 (n_6_2813), .C2 (n_6_1_973));
NAND2_X1 slo__sro_c30991 (.ZN (slo__sro_n27582), .A1 (slo__sro_n27583), .A2 (slo__sro_n27584));
INV_X1 slo__sro_c30975 (.ZN (slo__sro_n27573), .A (slo__sro_n8834));
NAND2_X1 slo__sro_c30976 (.ZN (slo__sro_n27572), .A1 (n_6_731), .A2 (n_6_1_729));
NAND2_X1 slo__sro_c30727 (.ZN (slo__sro_n27339), .A1 (opt_ipo_n45138), .A2 (n_6_1_448));
NAND2_X1 CLOCK_slo__sro_c58791 (.ZN (CLOCK_slo__sro_n53572), .A1 (slo__n28104), .A2 (n_6_1_238));
NAND2_X1 slo__sro_c30977 (.ZN (slo__sro_n27571), .A1 (slo__sro_n27572), .A2 (slo__sro_n27573));
AOI21_X2 slo__sro_c30978 (.ZN (n_6_1_723), .A (slo__sro_n27571), .B1 (n_6_763), .B2 (n_6_1_730));
NAND2_X1 CLOCK_sgo__sro_c51634 (.ZN (CLOCK_sgo__sro_n47370), .A1 (n_6_1602), .A2 (slo___n23215));
AOI21_X2 slo__sro_c31105 (.ZN (slo__sro_n27689), .A (slo__sro_n27690), .B1 (n_6_762), .B2 (n_6_1_730));
CLKBUF_X2 spw__c75857 (.Z (n_6_1_604), .A (spw__n67656));
NAND2_X1 slo__sro_c31140 (.ZN (slo__sro_n27728), .A1 (n_6_2198), .A2 (n_6_1_273));
AOI222_X2 CLOCK_slo__sro_c58576 (.ZN (n_6_1_632), .A1 (n_6_870), .A2 (n_6_1_660), .B1 (n_6_838)
    , .B2 (slo___n23463), .C1 (n_6_2517), .C2 (n_6_1_658));
AOI21_X2 CLOCK_slo__sro_c60699 (.ZN (CLOCK_slo__sro_n55168), .A (CLOCK_slo__sro_n55169)
    , .B1 (n_6_827), .B2 (n_6_1_695));
NOR2_X2 CLOCK_slo__sro_c61637 (.ZN (slo__sro_n37482), .A1 (slo__sro_n37483), .A2 (CLOCK_slo__sro_n55959));
NAND2_X1 slo__sro_c31397 (.ZN (slo__sro_n27973), .A1 (n_6_969), .A2 (slo___n23232));
NAND2_X1 slo__sro_c31306 (.ZN (slo__sro_n27893), .A1 (n_6_1_798), .A2 (n_6_2651));
NAND2_X1 slo__sro_c31307 (.ZN (slo__sro_n27892), .A1 (n_6_624), .A2 (n_6_1_800));
NAND2_X1 slo__sro_c31308 (.ZN (slo__sro_n27891), .A1 (slo__sro_n27892), .A2 (slo__sro_n27893));
AOI21_X2 slo__sro_c31309 (.ZN (CLOCK_slo__n50956), .A (slo__sro_n27891), .B1 (n_6_592), .B2 (n_6_1_799));
AND2_X1 slo__sro_c31237 (.ZN (slo__sro_n27823), .A1 (n_6_2411), .A2 (n_6_1_518));
AOI221_X2 slo__sro_c31238 (.ZN (slo__sro_n27822), .A (slo__sro_n27823), .B1 (n_6_1112)
    , .B2 (slo___n23277), .C1 (n_6_1144), .C2 (slo___n23268));
NAND2_X1 slo__sro_c31435 (.ZN (slo__sro_n28007), .A1 (n_6_817), .A2 (n_6_1_695));
NAND2_X1 slo__sro_c31436 (.ZN (slo__sro_n28006), .A1 (slo__sro_n28007), .A2 (slo__sro_n28008));
AOI21_X2 slo__sro_c31437 (.ZN (slo__sro_n7852), .A (slo__sro_n28006), .B1 (n_6_785), .B2 (n_6_1_694));
NAND2_X1 slo__sro_c31396 (.ZN (slo__sro_n27974), .A1 (opt_ipo_n25394), .A2 (n_6_1_588));
INV_X1 slo__L1_c1_c31503 (.ZN (slo__n28070), .A (slo__n28071));
INV_X2 slo__L1_c1_c31537 (.ZN (slo__n28104), .A (slo__n28105));
NAND2_X1 slo__sro_c31615 (.ZN (slo__sro_n28183), .A1 (n_6_2639), .A2 (n_6_1_798));
NAND2_X1 slo__sro_c31616 (.ZN (slo__sro_n28182), .A1 (n_6_612), .A2 (n_6_1_800));
NAND2_X1 slo__sro_c31617 (.ZN (slo__sro_n28181), .A1 (slo__sro_n28182), .A2 (slo__sro_n28183));
AOI21_X2 slo__sro_c31732 (.ZN (slo__sro_n28283), .A (slo__sro_n28284), .B1 (n_6_1531), .B2 (slo___n23247));
AOI21_X2 slo__sro_c31618 (.ZN (n_6_1_770), .A (slo__sro_n28181), .B1 (n_6_580), .B2 (n_6_1_799));
AND2_X1 slo__sro_c31780 (.ZN (slo__sro_n28334), .A1 (n_6_2379), .A2 (n_6_1_483));
AOI221_X2 slo__sro_c31781 (.ZN (slo__sro_n28333), .A (slo__sro_n28334), .B1 (n_6_1175)
    , .B2 (slo___n23364), .C1 (n_6_1207), .C2 (slo___n23466));
NAND2_X4 slo__sro_c31976 (.ZN (slo__sro_n28524), .A1 (slo__sro_n28525), .A2 (slo__sro_n28526));
AOI21_X4 slo__sro_c31871 (.ZN (slo__sro_n28419), .A (slo__sro_n28420), .B1 (n_6_1000), .B2 (slo___n23218));
AOI21_X1 slo__sro_c31977 (.ZN (slo__sro_n28523), .A (slo__sro_n28524), .B1 (n_6_748), .B2 (n_6_1_730));
NAND2_X1 CLOCK_sgo__sro_c51635 (.ZN (CLOCK_sgo__sro_n47369), .A1 (CLOCK_sgo__sro_n47370), .A2 (CLOCK_sgo__sro_n47371));
AND2_X1 slo__sro_c32043 (.ZN (slo__sro_n28592), .A1 (n_6_2494), .A2 (n_6_1_623));
NAND2_X1 slo__sro_c31729 (.ZN (slo__sro_n28286), .A1 (n_6_1_308), .A2 (n_6_2228));
NAND2_X1 slo__sro_c31730 (.ZN (slo__sro_n28285), .A1 (n_6_1499), .A2 (n_6_1_309));
INV_X1 slo__L1_c1_c31990 (.ZN (slo__n28538), .A (slo__n28539));
NAND2_X1 slo__sro_c31731 (.ZN (slo__sro_n28284), .A1 (slo__sro_n28285), .A2 (slo__sro_n28286));
NAND2_X1 CLOCK_sgo__sro_c51984 (.ZN (CLOCK_sgo__sro_n47663), .A1 (CLOCK_sgo__sro_n47664), .A2 (CLOCK_sgo__sro_n47665));
NAND2_X1 slo__sro_c32463 (.ZN (slo__sro_n28990), .A1 (n_6_2126), .A2 (n_6_1_203));
NAND2_X1 slo__sro_c32113 (.ZN (slo__sro_n28660), .A1 (n_6_2220), .A2 (n_6_1_308));
INV_X1 slo__sro_c32114 (.ZN (slo__sro_n28659), .A (slo__sro_n28660));
AOI221_X2 slo__sro_c32115 (.ZN (n_6_1_295), .A (slo__sro_n28659), .B1 (n_6_1491), .B2 (n_6_1_309)
    , .C1 (n_6_1523), .C2 (slo___n23247));
INV_X2 opt_ipo_c27440 (.ZN (opt_ipo_n24063), .A (slo__sro_n11594));
AOI221_X2 slo__sro_c32503 (.ZN (slo__sro_n29017), .A (slo__sro_n29018), .B1 (n_6_1795)
    , .B2 (n_6_1_134), .C1 (n_6_1827), .C2 (slo___n23404));
AOI21_X2 slo__sro_c32240 (.ZN (slo__sro_n28774), .A (slo__sro_n28775), .B1 (n_6_660), .B2 (n_6_1_764));
INV_X1 slo__sro_c32464 (.ZN (slo__sro_n28989), .A (slo__sro_n28990));
AOI221_X2 slo__sro_c32465 (.ZN (slo__sro_n14501), .A (slo__sro_n28989), .B1 (n_6_1714)
    , .B2 (slo___n23407), .C1 (n_6_1682), .C2 (n_6_1_204));
INV_X2 opt_ipo_c27452 (.ZN (opt_ipo_n24075), .A (n_6_1_107));
NAND2_X1 slo__sro_c32501 (.ZN (slo__sro_n29019), .A1 (n_6_2049), .A2 (n_6_1_133));
AOI221_X2 CLOCK_slo__sro_c59991 (.ZN (n_6_1_288), .A (slo__sro_n22964), .B1 (n_6_1484)
    , .B2 (n_6_1_309), .C1 (n_6_1516), .C2 (slo___n23247));
INV_X1 slo__sro_c32723 (.ZN (slo__sro_n29227), .A (n_6_1_308));
AND2_X1 slo__sro_c32664 (.ZN (slo__sro_n29176), .A1 (n_6_1467), .A2 (n_6_1_345));
AOI21_X1 slo__sro_c32863 (.ZN (slo__sro_n29362), .A (slo__sro_n29363), .B1 (n_6_977), .B2 (slo___n23232));
NAND2_X1 slo__sro_c32861 (.ZN (slo__sro_n29364), .A1 (n_6_1009), .A2 (slo___n23218));
NAND2_X1 slo__sro_c32697 (.ZN (slo__sro_n29207), .A1 (n_6_2406), .A2 (n_6_1_518));
NAND2_X1 slo__sro_c32698 (.ZN (slo__sro_n29206), .A1 (n_6_1107), .A2 (slo___n23277));
NAND2_X1 slo__sro_c32699 (.ZN (slo__sro_n29205), .A1 (slo__sro_n29206), .A2 (slo__sro_n29207));
NOR2_X2 slo__sro_c32665 (.ZN (slo__sro_n19751), .A1 (slo__sro_n19752), .A2 (slo__sro_n29176));
AOI21_X1 slo__sro_c32700 (.ZN (n_6_1_505), .A (slo__sro_n29205), .B1 (n_6_1139), .B2 (slo___n23268));
AOI21_X2 CLOCK_sgo__sro_c51636 (.ZN (n_6_1_208), .A (CLOCK_sgo__sro_n47369), .B1 (n_6_1634), .B2 (drc_ipo_n26601));
NOR2_X1 slo__sro_c32944 (.ZN (slo__sro_n29443), .A1 (slo__sro_n13738), .A2 (slo__sro_n29444));
AND2_X1 CLOCK_slo__sro_c56213 (.ZN (CLOCK_slo__sro_n51388), .A1 (n_6_1781), .A2 (CLOCK_sgo__n48020));
NAND2_X1 slo__sro_c33168 (.ZN (slo__sro_n29651), .A1 (slo__sro_n29653), .A2 (slo__sro_n29652));
NAND2_X1 slo__sro_c33166 (.ZN (slo__sro_n29653), .A1 (n_6_2299), .A2 (n_6_1_413));
NAND2_X1 slo__sro_c33192 (.ZN (slo__sro_n29675), .A1 (slo__sro_n29676), .A2 (slo__sro_n29677));
INV_X1 slo__sro_c32990 (.ZN (slo__sro_n29491), .A (slo__sro_n10518));
NAND2_X1 slo__sro_c32991 (.ZN (slo__sro_n29490), .A1 (n_6_1_869), .A2 (n_6_476));
NAND2_X1 slo__sro_c32992 (.ZN (slo__sro_n29489), .A1 (slo__sro_n29490), .A2 (slo__sro_n29491));
NAND2_X1 CLOCK_slo__sro_c61762 (.ZN (CLOCK_slo__sro_n56060), .A1 (CLOCK_sgo__n46950), .A2 (slo___n7881));
AND2_X2 CLOCK_slo__sro_c55615 (.ZN (CLOCK_slo__sro_n50850), .A1 (n_6_1507), .A2 (slo___n23247));
NAND2_X1 slo__sro_c33028 (.ZN (slo__sro_n29526), .A1 (CLOCK_sgo__n46945), .A2 (n_6_2872));
NAND2_X1 slo__sro_c33029 (.ZN (slo__sro_n29525), .A1 (n_6_180), .A2 (n_6_1_1045));
NAND2_X1 slo__sro_c33030 (.ZN (slo__sro_n29524), .A1 (slo__sro_n29525), .A2 (slo__sro_n29526));
AOI21_X1 slo__sro_c33031 (.ZN (slo__sro_n29523), .A (slo__sro_n29524), .B1 (n_6_148), .B2 (n_6_1_1044));
BUF_X4 CLOCK_sgo__L1_c1_c51020 (.Z (CLOCK_sgo__n46725), .A (Multiplier_19_PP_2));
NAND2_X1 slo__sro_c33340 (.ZN (slo__sro_n29824), .A1 (n_6_2745), .A2 (CLOCK_sgo__n46934));
NAND2_X1 slo__sro_c33289 (.ZN (slo__sro_n29774), .A1 (n_6_2672), .A2 (CLOCK_sgo__n46922));
INV_X1 slo__sro_c33290 (.ZN (slo__sro_n29773), .A (slo__sro_n29774));
INV_X1 slo__sro_c41784 (.ZN (slo__sro_n37843), .A (slo__sro_n30145));
NAND2_X1 slo__sro_c33341 (.ZN (slo__sro_n29823), .A1 (n_6_1_905), .A2 (n_6_433));
NAND2_X1 slo__sro_c33342 (.ZN (slo__sro_n29822), .A1 (slo__sro_n29823), .A2 (slo__sro_n29824));
AOI21_X1 slo__sro_c33343 (.ZN (n_6_1_888), .A (slo__sro_n29822), .B1 (n_6_401), .B2 (n_6_1_904));
NAND2_X2 slo__sro_c33381 (.ZN (slo__sro_n29858), .A1 (slo__sro_n29859), .A2 (slo__sro_n29860));
AOI21_X2 slo__sro_c33382 (.ZN (slo__sro_n29857), .A (slo__sro_n29858), .B1 (n_6_1719), .B2 (slo___n23407));
INV_X4 opt_ipo_c49450 (.ZN (opt_ipo_n45107), .A (n_6_1_125));
INV_X1 opt_ipo_c27543 (.ZN (opt_ipo_n24166), .A (slo__sro_n12865));
AOI21_X2 slo__sro_c33405 (.ZN (slo__sro_n4750), .A (slo__sro_n29880), .B1 (n_6_450), .B2 (n_6_1_869));
INV_X1 slo__sro_c33444 (.ZN (slo__sro_n29918), .A (slo__sro_n29919));
BUF_X4 spw__c75741 (.Z (n_6_1_107), .A (spw__n67541));
INV_X2 opt_ipo_c27550 (.ZN (opt_ipo_n24173), .A (n_6_1_880));
NAND2_X1 slo__sro_c33546 (.ZN (slo__sro_n30018), .A1 (slo__sro_n30019), .A2 (slo__sro_n30020));
AOI21_X1 slo__sro_c33547 (.ZN (slo__sro_n30017), .A (slo__sro_n30018), .B1 (n_6_784), .B2 (n_6_1_694));
NAND2_X1 slo__sro_c33560 (.ZN (slo__sro_n30032), .A1 (slo__sro_n30033), .A2 (slo__sro_n30034));
AOI21_X1 slo__sro_c33561 (.ZN (slo__sro_n30031), .A (slo__sro_n30032), .B1 (n_6_533), .B2 (n_6_1_834));
NAND2_X1 slo__sro_c33646 (.ZN (slo__sro_n30113), .A1 (n_6_2110), .A2 (n_6_1_203));
NAND2_X2 slo__sro_c33647 (.ZN (slo__sro_n30112), .A1 (n_6_1666), .A2 (n_6_1_204));
INV_X1 opt_ipo_c27567 (.ZN (opt_ipo_n24190), .A (slo__sro_n31654));
INV_X1 slo__sro_c33681 (.ZN (slo__sro_n30147), .A (n_6_2751));
NAND2_X1 slo__sro_c33599 (.ZN (slo__sro_n30073), .A1 (n_6_1_868), .A2 (n_6_2712));
BUF_X1 opt_ipo_c27573 (.Z (opt_ipo_n24196), .A (n_6_2027));
NAND2_X1 slo__sro_c33600 (.ZN (slo__sro_n30072), .A1 (n_6_495), .A2 (n_6_1_870));
NAND2_X1 slo__sro_c33601 (.ZN (slo__sro_n30071), .A1 (slo__sro_n30072), .A2 (slo__sro_n30073));
AOI21_X2 slo__sro_c33602 (.ZN (n_6_1_851), .A (slo__sro_n30071), .B1 (n_6_463), .B2 (n_6_1_869));
AOI21_X4 slo__sro_c33649 (.ZN (slo__sro_n30110), .A (slo__sro_n30111), .B1 (n_6_1698), .B2 (slo___n23407));
NOR2_X1 slo__sro_c33683 (.ZN (slo__sro_n30145), .A1 (slo__sro_n30147), .A2 (slo__sro_n30146));
INV_X4 slo__c42246 (.ZN (slo__n38218), .A (slo__sro_n15079));
NAND2_X1 slo__sro_c33747 (.ZN (slo__sro_n30209), .A1 (hfn_ipo_n30), .A2 (slo__n30589));
NAND2_X1 slo__sro_c33748 (.ZN (slo__sro_n30208), .A1 (Multiplicand[1]), .A2 (n_6_2913));
NAND2_X1 slo__sro_c33749 (.ZN (slo__sro_n30207), .A1 (slo__sro_n30208), .A2 (slo__sro_n30209));
AOI21_X1 slo__sro_c33750 (.ZN (n_6_1_1111), .A (slo__sro_n30207), .B1 (n_6_61), .B2 (n_6_1_1114));
NAND2_X1 slo__sro_c33809 (.ZN (slo__sro_n30265), .A1 (n_6_269), .A2 (n_6_1_974));
NAND2_X1 slo__sro_c33810 (.ZN (slo__sro_n30264), .A1 (slo__sro_n30265), .A2 (slo__sro_n30266));
AOI21_X1 slo__sro_c33811 (.ZN (slo__sro_n11034), .A (slo__sro_n30264), .B1 (n_6_301), .B2 (n_6_1_975));
NAND2_X2 slo__sro_c34967 (.ZN (slo__sro_n31361), .A1 (slo__sro_n31362), .A2 (slo__sro_n31363));
INV_X1 slo__sro_c33916 (.ZN (slo__sro_n30364), .A (slo__sro_n20420));
NAND2_X1 slo__sro_c33917 (.ZN (slo__sro_n30363), .A1 (n_6_852), .A2 (slo___n23463));
NAND2_X1 slo__sro_c33918 (.ZN (slo__sro_n30362), .A1 (slo__sro_n30363), .A2 (slo__sro_n30364));
AOI21_X2 slo__sro_c33919 (.ZN (n_6_1_646), .A (slo__sro_n30362), .B1 (n_6_884), .B2 (slo___n23451));
AOI21_X2 slo__sro_c34968 (.ZN (slo__sro_n4244), .A (slo__sro_n31361), .B1 (n_6_507), .B2 (n_6_1_870));
INV_X1 slo__sro_c34067 (.ZN (slo__sro_n30506), .A (slo__sro_n10378));
NAND2_X1 slo__sro_c34068 (.ZN (slo__sro_n30505), .A1 (n_6_411), .A2 (n_6_1_904));
INV_X2 opt_ipo_c27628 (.ZN (opt_ipo_n24251), .A (n_6_1_454));
AOI21_X2 slo__sro_c34070 (.ZN (n_6_1_898), .A (slo__sro_n30504), .B1 (n_6_443), .B2 (n_6_1_905));
NAND2_X2 slo__sro_c34287 (.ZN (slo__sro_n30705), .A1 (slo__sro_n30706), .A2 (slo__sro_n21212));
AOI21_X4 slo__sro_c34288 (.ZN (slo__sro_n30704), .A (slo__sro_n30705), .B1 (n_6_444), .B2 (n_6_1_905));
NAND2_X1 slo__sro_c34586 (.ZN (slo__sro_n30997), .A1 (n_6_1049), .A2 (n_6_1_554));
INV_X1 slo__sro_c34506 (.ZN (slo__sro_n30924), .A (n_6_2116));
INV_X1 slo__sro_c34507 (.ZN (slo__sro_n30923), .A (n_6_1_203));
NOR2_X1 slo__sro_c34508 (.ZN (slo__sro_n30922), .A1 (slo__sro_n30924), .A2 (slo__sro_n30923));
NAND2_X2 CLOCK_slo__sro_c58456 (.ZN (CLOCK_slo__sro_n53277), .A1 (CLOCK_slo__sro_n53278), .A2 (slo__sro_n27728));
NAND2_X2 slo__sro_c34587 (.ZN (slo__sro_n30996), .A1 (slo__sro_n30997), .A2 (slo__sro_n30998));
AOI21_X4 slo__sro_c34588 (.ZN (slo__sro_n30995), .A (slo__sro_n30996), .B1 (n_6_1081), .B2 (slo___n23457));
AOI21_X2 slo__sro_c34644 (.ZN (slo__sro_n31050), .A (slo__sro_n31051), .B1 (n_6_1330), .B2 (slo___n43257));
INV_X1 slo__sro_c34679 (.ZN (slo__sro_n31088), .A (slo__sro_n31089));
AOI221_X2 slo__sro_c34680 (.ZN (slo__sro_n31087), .A (slo__sro_n31088), .B1 (n_6_1092)
    , .B2 (slo___n23277), .C1 (n_6_1124), .C2 (slo___n23268));
NAND2_X1 slo__sro_c34813 (.ZN (slo__sro_n31218), .A1 (slo__sro_n31219), .A2 (slo__sro_n31220));
INV_X4 opt_ipo_c27662 (.ZN (opt_ipo_n24285), .A (slo__sro_n37401));
AOI21_X2 slo__sro_c34814 (.ZN (n_6_1_479), .A (slo__sro_n31218), .B1 (n_6_1212), .B2 (slo___n23466));
NAND2_X1 slo__sro_c34832 (.ZN (slo__sro_n31236), .A1 (n_6_1289), .A2 (n_6_1_414));
NAND2_X1 slo__sro_c34833 (.ZN (slo__sro_n31235), .A1 (slo__sro_n31236), .A2 (slo__sro_n31237));
AOI21_X1 slo__sro_c34834 (.ZN (slo__sro_n31234), .A (slo__sro_n31235), .B1 (n_6_1321), .B2 (slo___n43257));
NAND2_X1 slo__sro_c35181 (.ZN (slo__sro_n31560), .A1 (slo__sro_n31561), .A2 (slo__sro_n31562));
CLKBUF_X2 CLOCK_opt_ipo_c50085 (.Z (CLOCK_opt_ipo_n45742), .A (CLOCK_opt_ipo_n45744));
NAND2_X2 slo__sro_c34904 (.ZN (slo__sro_n31307), .A1 (n_6_483), .A2 (n_6_1_870));
NAND2_X2 slo__sro_c34905 (.ZN (slo__sro_n31306), .A1 (slo__sro_n31307), .A2 (slo__sro_n11071));
AOI21_X2 slo__sro_c34906 (.ZN (n_6_1_839), .A (slo__sro_n31306), .B1 (n_6_451), .B2 (n_6_1_869));
NAND2_X1 CLOCK_sgo__sro_c51500 (.ZN (CLOCK_sgo__sro_n47263), .A1 (n_6_1_273), .A2 (slo___n17633));
NAND2_X1 slo__sro_c35097 (.ZN (slo__sro_n31484), .A1 (n_6_617), .A2 (n_6_1_800));
INV_X1 slo__sro_c34965 (.ZN (slo__sro_n31363), .A (slo__sro_n4245));
NAND2_X1 slo__sro_c34966 (.ZN (slo__sro_n31362), .A1 (n_6_1_869), .A2 (n_6_475));
NAND2_X1 slo__sro_c35098 (.ZN (slo__sro_n31483), .A1 (slo__sro_n16242), .A2 (slo__sro_n31484));
AOI21_X2 slo__sro_c35099 (.ZN (n_6_1_775), .A (slo__sro_n31483), .B1 (n_6_585), .B2 (n_6_1_799));
AOI21_X2 slo__sro_c35182 (.ZN (slo__sro_n31559), .A (slo__sro_n31560), .B1 (n_6_903), .B2 (slo___n23367));
INV_X1 slo__sro_c35272 (.ZN (slo__sro_n31646), .A (slo__sro_n18863));
INV_X1 opt_ipo_c27703 (.ZN (opt_ipo_n24326), .A (slo__sro_n27836));
NAND2_X2 slo__sro_c35274 (.ZN (slo__sro_n31644), .A1 (slo__sro_n31645), .A2 (slo__sro_n31646));
AOI21_X4 slo__sro_c35275 (.ZN (n_6_1_966), .A (slo__sro_n31644), .B1 (n_6_313), .B2 (n_6_1_975));
NAND2_X1 slo__sro_c35303 (.ZN (slo__sro_n31671), .A1 (n_6_284), .A2 (n_6_1_974));
NAND2_X1 slo__sro_c35304 (.ZN (slo__sro_n31670), .A1 (slo__sro_n31671), .A2 (slo__sro_n31672));
INV_X1 CLOCK_slo__sro_c60146 (.ZN (CLOCK_slo__sro_n54706), .A (CLOCK_slo__sro_n54707));
NAND2_X1 slo__sro_c35455 (.ZN (slo__sro_n31819), .A1 (CLOCK_opt_ipo_n45873), .A2 (CLOCK_sgo__n46934));
NAND2_X1 slo__sro_c35437 (.ZN (slo__sro_n31801), .A1 (n_6_2438), .A2 (n_6_1_553));
NAND2_X1 slo__sro_c35438 (.ZN (slo__sro_n31800), .A1 (n_6_1044), .A2 (n_6_1_554));
NAND2_X1 slo__sro_c35439 (.ZN (slo__sro_n31799), .A1 (slo__sro_n31800), .A2 (slo__sro_n31801));
AOI21_X2 slo__sro_c35440 (.ZN (slo__sro_n31798), .A (slo__sro_n31799), .B1 (n_6_1076), .B2 (slo___n23457));
NAND2_X1 slo__sro_c35457 (.ZN (slo__sro_n31817), .A1 (slo__sro_n31818), .A2 (slo__sro_n31819));
AOI21_X2 slo__sro_c35458 (.ZN (slo__sro_n31816), .A (slo__sro_n31817), .B1 (n_6_421), .B2 (n_6_1_905));
BUF_X4 opt_ipo_c27735 (.Z (opt_ipo_n24358), .A (sgo__n691));
AOI21_X2 slo__sro_c35681 (.ZN (slo__sro_n32026), .A (slo__sro_n32027), .B1 (n_6_584), .B2 (n_6_1_799));
NAND2_X2 slo__mro_c35505 (.ZN (slo__sro_n22554), .A1 (n_6_344), .A2 (n_6_1_939));
NAND2_X1 slo__sro_c35678 (.ZN (slo__sro_n32029), .A1 (slo___n15116), .A2 (n_6_1_798));
NAND2_X1 slo__sro_c35679 (.ZN (slo__sro_n32028), .A1 (n_6_616), .A2 (n_6_1_800));
NAND2_X2 slo__sro_c35698 (.ZN (slo__sro_n32045), .A1 (slo__sro_n32046), .A2 (slo__sro_n7371));
AOI21_X4 slo__sro_c35699 (.ZN (slo__sro_n32044), .A (slo__sro_n32045), .B1 (n_6_899), .B2 (slo___n23367));
INV_X1 slo__sro_c35774 (.ZN (slo__sro_n32119), .A (n_6_1_518));
NOR2_X1 slo__sro_c35775 (.ZN (slo__sro_n32118), .A1 (slo__sro_n32120), .A2 (slo__sro_n32119));
AOI221_X2 slo__sro_c35776 (.ZN (slo__sro_n32117), .A (slo__sro_n32118), .B1 (n_6_1125)
    , .B2 (slo___n23268), .C1 (n_6_1093), .C2 (slo___n23277));
NAND2_X1 CLOCK_slo__sro_c69872 (.ZN (CLOCK_slo__sro_n62931), .A1 (n_6_917), .A2 (slo___n23367));
NAND2_X1 CLOCK_slo__sro_c53264 (.ZN (CLOCK_slo__sro_n48741), .A1 (n_6_1607), .A2 (slo___n23215));
NAND2_X1 slo__sro_c35838 (.ZN (slo__sro_n32185), .A1 (slo__n13799), .A2 (n_6_2895));
INV_X1 slo__sro_c35819 (.ZN (slo__sro_n32166), .A (slo__sro_n20666));
NAND2_X1 slo__sro_c35820 (.ZN (slo__sro_n32165), .A1 (slo___n23215), .A2 (n_6_1628));
NAND2_X1 slo__sro_c35821 (.ZN (slo__sro_n32164), .A1 (slo__sro_n32165), .A2 (slo__sro_n32166));
AOI21_X2 slo__sro_c35822 (.ZN (slo__sro_n32163), .A (slo__sro_n32164), .B1 (n_6_1660), .B2 (drc_ipo_n26601));
NAND2_X1 slo__sro_c35839 (.ZN (slo__sro_n32184), .A1 (n_6_1_1080), .A2 (n_6_108));
NAND2_X1 slo__sro_c35840 (.ZN (slo__sro_n32183), .A1 (slo__sro_n32184), .A2 (slo__sro_n32185));
AOI21_X1 slo__sro_c35841 (.ZN (slo__sro_n32182), .A (slo__sro_n32183), .B1 (n_6_76), .B2 (n_6_1_1079));
NAND2_X2 slo__sro_c35860 (.ZN (slo__sro_n32202), .A1 (slo__sro_n32203), .A2 (slo__sro_n32204));
AOI21_X4 slo__sro_c35861 (.ZN (n_6_1_162), .A (slo__sro_n32202), .B1 (n_6_1786), .B2 (CLOCK_sgo__n48020));
NAND2_X1 slo__sro_c35980 (.ZN (slo__sro_n32318), .A1 (n_6_1542), .A2 (n_6_1_274));
NAND2_X1 slo__sro_c36147 (.ZN (slo__sro_n32472), .A1 (n_6_1475), .A2 (n_6_1_309));
NAND2_X1 slo__sro_c35981 (.ZN (slo__sro_n32317), .A1 (slo__sro_n32318), .A2 (slo__sro_n32319));
AOI21_X2 slo__sro_c35982 (.ZN (slo__sro_n32316), .A (slo__sro_n32317), .B1 (n_6_1574), .B2 (slo___n23244));
AND2_X1 slo__sro_c36022 (.ZN (slo__sro_n32358), .A1 (n_6_2867), .A2 (CLOCK_sgo__n46945));
AOI221_X1 slo__sro_c36023 (.ZN (slo__sro_n32357), .A (slo__sro_n32358), .B1 (n_6_175)
    , .B2 (n_6_1_1045), .C1 (n_6_143), .C2 (n_6_1_1044));
AOI21_X2 CLOCK_slo__sro_c69874 (.ZN (slo__sro_n19727), .A (CLOCK_slo__sro_n62930)
    , .B1 (n_6_949), .B2 (n_6_1_625));
INV_X2 opt_ipo_c27808 (.ZN (opt_ipo_n24431), .A (CLOCK_slo__sro_n53196));
NAND2_X2 slo__sro_c36148 (.ZN (slo__sro_n32471), .A1 (slo__sro_n32472), .A2 (slo__sro_n32473));
INV_X2 opt_ipo_c49481 (.ZN (opt_ipo_n45138), .A (CLOCK_slo__sro_n52124));
NAND2_X1 slo__mro_c36209 (.ZN (slo__mro_n32529), .A1 (n_6_1736), .A2 (n_6_1_169));
AOI221_X2 slo__sro_c36414 (.ZN (slo__sro_n32716), .A (slo__sro_n32717), .B1 (n_6_811)
    , .B2 (n_6_1_695), .C1 (n_6_779), .C2 (n_6_1_694));
AOI21_X4 slo__mro_c36956 (.ZN (slo__mro_n33299), .A (slo__mro_n33302), .B1 (slo__mro_n33301), .B2 (slo__mro_n33300));
OAI21_X1 slo__mro_c36719 (.ZN (slo__sro_n11216), .A (slo__sro_n11218), .B1 (opt_ipo_n45556), .B2 (slo__mro_n33047));
NAND2_X1 slo__sro_c38247 (.ZN (slo__sro_n34607), .A1 (slo__sro_n34608), .A2 (slo__sro_n34609));
AND2_X1 slo__sro_c37195 (.ZN (slo__sro_n33527), .A1 (n_6_2192), .A2 (n_6_1_273));
AOI221_X2 slo__sro_c37196 (.ZN (slo__sro_n33526), .A (slo__sro_n33527), .B1 (n_6_1558)
    , .B2 (n_6_1_274), .C1 (n_6_1590), .C2 (slo___n23244));
AOI222_X2 slo__sro_c37030 (.ZN (slo__sro_n33373), .A1 (n_6_1334), .A2 (slo___n43257)
    , .B1 (n_6_1302), .B2 (n_6_1_414), .C1 (CLOCK_slo__n57799), .C2 (n_6_1_413));
AOI21_X2 slo__sro_c37270 (.ZN (slo__sro_n33595), .A (slo__sro_n33596), .B1 (n_6_1720), .B2 (slo___n23407));
AOI222_X1 slo__sro_c37708 (.ZN (slo__sro_n34095), .A1 (n_6_843), .A2 (slo___n23463)
    , .B1 (n_6_875), .B2 (n_6_1_660), .C1 (slo___n17357), .C2 (n_6_1_658));
NAND2_X2 slo__sro_c38399 (.ZN (slo__sro_n34756), .A1 (slo__sro_n34757), .A2 (slo__sro_n34758));
INV_X1 slo__sro_c37861 (.ZN (slo__sro_n34247), .A (slo__sro_n34248));
INV_X1 CLOCK_slo__c61256 (.ZN (CLOCK_slo__n55658), .A (slo__sro_n19567));
NAND2_X1 CLOCK_slo__sro_c56905 (.ZN (CLOCK_slo__sro_n51959), .A1 (n_6_332), .A2 (n_6_1_939));
AOI222_X2 slo__sro_c37352 (.ZN (slo__sro_n33677), .A1 (n_6_128), .A2 (n_6_1_1044)
    , .B1 (n_6_160), .B2 (n_6_1_1045), .C1 (n_6_2852), .C2 (CLOCK_sgo__n46945));
AOI221_X2 slo__sro_c38592 (.ZN (CLOCK_slo__n48588), .A (slo__sro_n34941), .B1 (n_6_294)
    , .B2 (n_6_1_975), .C1 (n_6_262), .C2 (n_6_1_974));
INV_X1 slo__sro_c37468 (.ZN (slo__sro_n33789), .A (slo__sro_n33790));
NAND2_X1 CLOCK_slo__sro_c55424 (.ZN (CLOCK_slo__sro_n50682), .A1 (n_6_2500), .A2 (n_6_1_623));
INV_X1 slo__mro_c36882 (.ZN (slo__mro_n33239), .A (n_6_1683));
INV_X1 slo__mro_c36883 (.ZN (slo__mro_n33238), .A (n_6_1_204));
AOI221_X2 slo__sro_c38262 (.ZN (slo__sro_n34620), .A (slo__sro_n34621), .B1 (n_6_788)
    , .B2 (n_6_1_694), .C1 (n_6_820), .C2 (n_6_1_695));
NAND2_X2 slo__sro_c38398 (.ZN (slo__sro_n34757), .A1 (n_6_1479), .A2 (n_6_1_309));
AOI221_X2 slo__sro_c38855 (.ZN (slo__sro_n35197), .A (slo__sro_n35198), .B1 (n_6_198)
    , .B2 (n_6_1_1009), .C1 (n_6_230), .C2 (n_6_1_1010));
NAND2_X1 slo__sro_c38795 (.ZN (slo__sro_n35145), .A1 (n_6_2165), .A2 (n_6_1_238));
AND2_X1 slo__sro_c38192 (.ZN (slo__sro_n34554), .A1 (n_6_2195), .A2 (n_6_1_273));
INV_X1 opt_ipo_c27880 (.ZN (opt_ipo_n24503), .A (n_6_1_993));
AOI21_X1 slo__mro_c36919 (.ZN (slo__mro_n33267), .A (n_6_1_62), .B1 (n_6_1949), .B2 (n_6_1_64));
NAND2_X1 slo__mro_c36678 (.ZN (slo__mro_n33015), .A1 (n_6_360), .A2 (n_6_1_940));
NAND2_X1 slo__mro_c36679 (.ZN (slo__mro_n33014), .A1 (slo__mro_n33015), .A2 (slo__sro_n22350));
INV_X1 slo__sro_c39053 (.ZN (slo__sro_n35378), .A (slo__sro_n13545));
NAND2_X1 slo__sro_c39054 (.ZN (slo__sro_n35377), .A1 (n_6_1_905), .A2 (n_6_434));
BUF_X4 CLOCK_sgo__L2_c2_c51051 (.Z (CLOCK_sgo__n46808), .A (drc_ipoPP_3PP_0));
NAND2_X1 slo__sro_c38984 (.ZN (slo__sro_n35312), .A1 (slo__sro_n35313), .A2 (slo__sro_n4661));
AND2_X1 slo__sro_c38912 (.ZN (slo__sro_n35250), .A1 (n_6_2610), .A2 (n_6_1_763));
INV_X1 CLOCK_sgo__sro_c51835 (.ZN (CLOCK_sgo__sro_n47541), .A (n_6_1800));
AOI21_X2 slo__sro_c38842 (.ZN (slo__sro_n35183), .A (slo__sro_n35184), .B1 (n_6_693), .B2 (n_6_1_765));
AOI222_X2 slo__sro_c38868 (.ZN (n_6_1_329), .A1 (n_6_1458), .A2 (n_6_1_345), .B1 (n_6_1426)
    , .B2 (slo___n23229), .C1 (n_6_2250), .C2 (n_6_1_343));
INV_X1 CLOCK_slo__c72160 (.ZN (CLOCK_slo__n64837), .A (slo__sro_n31654));
INV_X2 slo__L1_c1_c38767 (.ZN (slo__n35114), .A (slo__n35115));
NAND2_X2 CLOCK_slo__sro_c53835 (.ZN (CLOCK_slo__sro_n49243), .A1 (n_6_1113), .A2 (slo___n23277));
INV_X2 opt_ipo_c27918 (.ZN (opt_ipo_n24541), .A (n_6_1_217));
AOI21_X2 slo__sro_c38248 (.ZN (slo__sro_n34606), .A (slo__sro_n34607), .B1 (n_6_442), .B2 (n_6_1_905));
AND2_X1 slo__sro_c38591 (.ZN (slo__sro_n34941), .A1 (n_6_2796), .A2 (n_6_1_973));
AND2_X1 slo__sro_c37644 (.ZN (slo__sro_n34035), .A1 (n_6_1_782), .A2 (n_6_1_763));
INV_X2 CLOCK_slo__c64511 (.ZN (CLOCK_slo__n58182), .A (CLOCK_slo__sro_n50400));
NAND2_X1 slo__sro_c37860 (.ZN (slo__sro_n34248), .A1 (n_6_2857), .A2 (CLOCK_sgo__n46945));
NAND2_X1 slo__sro_c38841 (.ZN (slo__sro_n35184), .A1 (slo__sro_n35185), .A2 (slo__sro_n35186));
AOI21_X2 slo__sro_c38985 (.ZN (n_6_1_233), .A (slo__sro_n35312), .B1 (n_6_1659), .B2 (drc_ipo_n26601));
NAND2_X1 slo__sro_c39055 (.ZN (slo__sro_n35376), .A1 (slo__sro_n35377), .A2 (slo__sro_n35378));
AOI21_X1 slo__sro_c39056 (.ZN (slo__sro_n35375), .A (slo__sro_n35376), .B1 (n_6_402), .B2 (n_6_1_904));
AOI222_X2 slo__sro_c39023 (.ZN (n_6_1_1037), .A1 (n_6_186), .A2 (n_6_1_1045), .B1 (n_6_154)
    , .B2 (n_6_1_1044), .C1 (slo__sro_n23158), .C2 (CLOCK_sgo__n46945));
AND2_X1 slo__sro_c39096 (.ZN (slo__sro_n35419), .A1 (n_6_2709), .A2 (n_6_1_868));
NAND2_X1 CLOCK_slo__sro_c72470 (.ZN (CLOCK_slo__sro_n65090), .A1 (n_6_1_1010), .A2 (n_6_236));
INV_X1 slo__c40241 (.ZN (slo__n36492), .A (CLOCK_slo__sro_n56126));
INV_X1 slo__sro_c40466 (.ZN (slo__sro_n36683), .A (slo__sro_n36684));
AOI21_X2 CLOCK_slo__c72951 (.ZN (CLOCK_slo__n65456), .A (CLOCK_slo__sro_n53405), .B1 (n_6_1071), .B2 (slo___n23457));
NAND2_X2 slo__sro_c31975 (.ZN (slo__sro_n28525), .A1 (n_6_716), .A2 (n_6_1_729));
NAND2_X2 slo__sro_c31870 (.ZN (slo__sro_n28420), .A1 (slo__sro_n28421), .A2 (slo__sro_n28422));
AND2_X1 slo__sro_c40330 (.ZN (slo__sro_n36567), .A1 (n_6_2125), .A2 (n_6_1_203));
NAND2_X2 CLOCK_slo__c67591 (.ZN (slo__sro_n2968), .A1 (CLOCK_sgo__sro_n47846), .A2 (CLOCK_sgo__sro_n47847));
AOI221_X2 slo__sro_c39465 (.ZN (slo__sro_n15342), .A (slo__sro_n15343), .B1 (n_6_1651)
    , .B2 (drc_ipo_n26601), .C1 (n_6_1619), .C2 (slo___n23215));
NAND2_X1 slo__sro_c39378 (.ZN (slo__sro_n35684), .A1 (n_6_2894), .A2 (slo__n13799));
NAND2_X1 slo__sro_c39379 (.ZN (slo__sro_n35683), .A1 (n_6_107), .A2 (n_6_1_1080));
NAND2_X1 slo__sro_c39380 (.ZN (slo__sro_n35682), .A1 (slo__sro_n35684), .A2 (slo__sro_n35683));
NAND2_X1 CLOCK_slo__sro_c65215 (.ZN (CLOCK_slo__sro_n58766), .A1 (n_6_2375), .A2 (n_6_1_483));
NAND2_X1 CLOCK_slo__sro_c68172 (.ZN (CLOCK_slo__sro_n61396), .A1 (n_6_1333), .A2 (slo___n43257));
AOI21_X1 slo__sro_c39381 (.ZN (slo__sro_n35681), .A (slo__sro_n35682), .B1 (n_6_75), .B2 (n_6_1_1079));
AOI222_X2 slo__sro_c39804 (.ZN (slo__sro_n36088), .A1 (n_6_1424), .A2 (slo___n23229)
    , .B1 (n_6_1456), .B2 (n_6_1_345), .C1 (n_6_2248), .C2 (n_6_1_343));
AOI21_X1 slo__sro_c40640 (.ZN (n_6_1_514), .A (slo__sro_n36835), .B1 (n_6_1148), .B2 (slo___n23268));
AOI222_X2 slo__sro_c40824 (.ZN (n_6_1_396), .A1 (n_6_1295), .A2 (n_6_1_414), .B1 (n_6_1327)
    , .B2 (slo___n43257), .C1 (n_6_2309), .C2 (n_6_1_413));
NAND2_X1 slo__sro_c41084 (.ZN (slo__sro_n37224), .A1 (n_6_2911), .A2 (slo__n13799));
INV_X1 slo__sro_c40159 (.ZN (slo__sro_n36419), .A (n_6_2492));
NAND2_X1 slo__sro_c41085 (.ZN (slo__sro_n37223), .A1 (n_6_1_1079), .A2 (n_6_92));
AOI222_X2 slo__sro_c40728 (.ZN (slo__sro_n36913), .A1 (n_6_1096), .A2 (slo___n23277)
    , .B1 (n_6_1128), .B2 (slo___n23268), .C1 (n_6_2395), .C2 (n_6_1_518));
AOI221_X1 slo__sro_c40612 (.ZN (slo__sro_n36810), .A (n_6_1_552), .B1 (n_6_1086), .B2 (slo___n23457)
    , .C1 (n_6_1054), .C2 (n_6_1_554));
OR2_X4 slo__c40704 (.ZN (slo__sro_n23158), .A1 (slo__sro_n7833), .A2 (slo__sro_n23159));
AOI221_X2 slo__sro_c40537 (.ZN (n_6_1_574), .A (slo__sro_n9745), .B1 (n_6_978), .B2 (slo___n23232)
    , .C1 (n_6_1010), .C2 (slo___n23218));
AOI221_X2 slo__sro_c40467 (.ZN (n_6_1_650), .A (slo__sro_n36683), .B1 (n_6_888), .B2 (slo___n23451)
    , .C1 (n_6_856), .C2 (slo___n23463));
INV_X1 slo__sro_c39306 (.ZN (slo__sro_n35618), .A (slo__sro_n8171));
NAND2_X2 slo__sro_c39307 (.ZN (slo__sro_n35617), .A1 (n_6_355), .A2 (n_6_1_940));
NAND2_X1 CLOCK_slo__sro_c70256 (.ZN (CLOCK_slo__sro_n63269), .A1 (n_6_271), .A2 (n_6_1_974));
NAND2_X1 CLOCK_slo__sro_c60145 (.ZN (CLOCK_slo__sro_n54707), .A1 (n_6_2048), .A2 (n_6_1_133));
NAND2_X1 slo__sro_c41069 (.ZN (slo__sro_n37210), .A1 (n_6_665), .A2 (n_6_1_764));
NAND2_X1 CLOCK_slo__sro_c64675 (.ZN (CLOCK_slo__sro_n58315), .A1 (n_6_2638), .A2 (n_6_1_798));
INV_X1 slo__c40082 (.ZN (slo__n36345), .A (CLOCK_slo__sro_n52466));
INV_X2 slo__c39936 (.ZN (slo__n36214), .A (n_6_1_1085));
NAND2_X1 slo__sro_c40890 (.ZN (slo__sro_n37055), .A1 (n_6_176), .A2 (n_6_1_1045));
AOI21_X2 slo__sro_c40891 (.ZN (slo__sro_n37054), .A (slo__sro_n22874), .B1 (n_6_144), .B2 (n_6_1_1044));
AND2_X2 slo__sro_c40892 (.ZN (slo__sro_n37053), .A1 (slo__sro_n37054), .A2 (slo__sro_n37055));
NAND2_X1 slo__sro_c41189 (.ZN (slo__sro_n37306), .A1 (slo__sro_n37307), .A2 (slo__sro_n37308));
NAND2_X1 CLOCK_slo__sro_c66877 (.ZN (CLOCK_slo__sro_n60278), .A1 (n_6_2682), .A2 (CLOCK_sgo__n46922));
AOI21_X2 slo__sro_c41272 (.ZN (slo__sro_n37387), .A (slo__sro_n37388), .B1 (n_6_676), .B2 (n_6_1_765));
INV_X1 slo__sro_c41284 (.ZN (slo__sro_n37404), .A (n_6_802));
INV_X1 slo__sro_c41285 (.ZN (slo__sro_n37403), .A (n_6_1_695));
NAND2_X1 slo__sro_c41269 (.ZN (slo__sro_n37390), .A1 (n_6_1_763), .A2 (n_6_2608));
NAND2_X1 slo__sro_c41270 (.ZN (slo__sro_n37389), .A1 (n_6_1_764), .A2 (n_6_644));
OAI21_X2 slo__sro_c41286 (.ZN (slo__sro_n37402), .A (slo__sro_n37405), .B1 (slo__sro_n37404), .B2 (slo__sro_n37403));
AOI21_X4 slo__sro_c41287 (.ZN (slo__sro_n37401), .A (slo__sro_n37402), .B1 (n_6_770), .B2 (n_6_1_694));
NAND2_X1 slo__sro_c41385 (.ZN (slo__sro_n37483), .A1 (slo__sro_n37484), .A2 (slo__sro_n37485));
INV_X1 slo__c41300 (.ZN (slo__n37415), .A (slo__sro_n10270));
INV_X2 slo__c41328 (.ZN (slo__n37437), .A (slo__sro_n35163));
INV_X1 slo__c41361 (.ZN (slo__n37463), .A (n_6_1_779));
NAND2_X1 slo__sro_c41343 (.ZN (slo__sro_n37454), .A1 (CLOCK_sgo__n46950), .A2 (n_6_2849));
NAND2_X1 slo__sro_c41344 (.ZN (slo__sro_n37453), .A1 (n_6_1_1009), .A2 (n_6_220));
NAND2_X1 CLOCK_slo__sro_c54529 (.ZN (CLOCK_slo__sro_n49863), .A1 (slo__sro_n6090), .A2 (CLOCK_slo__sro_n49864));
BUF_X4 opt_ipo_c28075 (.Z (opt_ipo_n24698), .A (sgo__n1314));
NOR2_X2 CLOCK_slo__sro_c61697 (.ZN (n_6_1_1071), .A1 (slo__sro_n8430), .A2 (CLOCK_slo__sro_n56009));
AOI21_X1 slo__sro_c41456 (.ZN (slo__sro_n37540), .A (slo__sro_n29773), .B1 (n_6_550), .B2 (n_6_1_835));
INV_X4 slo__c41406 (.ZN (slo__n37502), .A (slo__sro_n40459));
INV_X2 opt_ipo_c28084 (.ZN (opt_ipo_n24707), .A (slo__sro_n14179));
NAND2_X1 slo__sro_c41785 (.ZN (slo__sro_n37842), .A1 (n_6_439), .A2 (n_6_1_905));
INV_X1 slo__c41468 (.ZN (slo__n37549), .A (n_6_1_879));
INV_X2 slo__c42001 (.ZN (slo__n38018), .A (n_6_1_470));
AOI222_X2 slo__sro_c41948 (.ZN (slo__sro_n37974), .A1 (n_6_1291), .A2 (n_6_1_414)
    , .B1 (n_6_1323), .B2 (slo___n43257), .C1 (n_6_2305), .C2 (n_6_1_413));
NAND2_X2 slo__sro_c41786 (.ZN (slo__sro_n37841), .A1 (slo__sro_n37842), .A2 (slo__sro_n37843));
INV_X1 opt_ipo_c28098 (.ZN (opt_ipo_n24721), .A (n_6_1_329));
NAND2_X1 slo__sro_c40222 (.ZN (slo__sro_n36479), .A1 (n_6_1_553), .A2 (n_6_2426));
INV_X4 opt_ipo_c28104 (.ZN (opt_ipo_n24727), .A (slo__sro_n19420));
AOI222_X2 slo__sro_c39758 (.ZN (slo__sro_n36045), .A1 (n_6_1677), .A2 (slo___n23239)
    , .B1 (n_6_1709), .B2 (slo___n23407), .C1 (n_6_2121), .C2 (n_6_1_203));
INV_X1 slo__c42785 (.ZN (slo__n38665), .A (n_6_1_1052));
INV_X1 slo__c42045 (.ZN (slo__n38056), .A (slo__sro_n15043));
INV_X2 slo__c42261 (.ZN (slo__n38227), .A (slo__sro_n5416));
INV_X1 slo__c42280 (.ZN (slo__n38240), .A (slo__sro_n29380));
INV_X2 opt_ipo_c28120 (.ZN (opt_ipo_n24743), .A (n_6_1_580));
NAND2_X2 CLOCK_slo__sro_c58616 (.ZN (CLOCK_slo__sro_n53419), .A1 (CLOCK_slo__sro_n53420), .A2 (slo__sro_n27339));
NAND2_X1 slo__sro_c42808 (.ZN (slo__sro_n38687), .A1 (n_6_2729), .A2 (CLOCK_sgo__n46934));
NAND2_X1 slo__sro_c42476 (.ZN (slo__sro_n38409), .A1 (slo__sro_n38410), .A2 (slo__sro_n38411));
NAND2_X1 CLOCK_slo__sro_c54883 (.ZN (CLOCK_slo__sro_n50188), .A1 (n_6_2514), .A2 (n_6_1_658));
NAND2_X1 slo__sro_c42809 (.ZN (slo__sro_n38686), .A1 (n_6_417), .A2 (n_6_1_905));
INV_X1 slo__sro_c42347 (.ZN (slo__sro_n38300), .A (opt_ipo_n45366));
INV_X1 slo__sro_c42348 (.ZN (slo__sro_n38299), .A (n_6_1_588));
NOR2_X1 slo__sro_c42349 (.ZN (slo__sro_n38298), .A1 (slo__sro_n38300), .A2 (slo__sro_n38299));
AOI221_X2 slo__sro_c42350 (.ZN (n_6_1_580), .A (slo__sro_n38298), .B1 (n_6_984), .B2 (slo___n23232)
    , .C1 (n_6_1016), .C2 (slo___n23218));
INV_X1 slo__c42770 (.ZN (slo__n38656), .A (slo__sro_n16180));
INV_X1 slo__c42662 (.ZN (slo__n38566), .A (n_6_1_882));
BUF_X16 slo__c42707 (.Z (slo__n38599), .A (sgo__n1311));
NAND2_X1 slo__sro_c42810 (.ZN (slo__sro_n38685), .A1 (slo__sro_n38686), .A2 (slo__sro_n38687));
AOI21_X1 slo__sro_c42811 (.ZN (slo__sro_n38684), .A (slo__sro_n38685), .B1 (n_6_385), .B2 (n_6_1_904));
NAND2_X1 CLOCK_sgo__sro_c51477 (.ZN (CLOCK_sgo__sro_n47245), .A1 (CLOCK_sgo__n48020), .A2 (n_6_1779));
AOI222_X2 slo__sro_c41759 (.ZN (slo__sro_n37819), .A1 (n_6_1002), .A2 (slo___n23218)
    , .B1 (n_6_970), .B2 (slo___n23232), .C1 (n_6_2459), .C2 (n_6_1_588));
INV_X2 opt_ipo_c28161 (.ZN (opt_ipo_n24784), .A (n_6_1_1069));
NAND2_X1 slo__sro_c42876 (.ZN (slo__sro_n38745), .A1 (slo__sro_n38746), .A2 (slo__sro_n38747));
AOI21_X1 slo__sro_c42877 (.ZN (slo__sro_n38744), .A (slo__sro_n38745), .B1 (n_6_880), .B2 (n_6_1_660));
NAND2_X1 slo__sro_c42889 (.ZN (slo__sro_n38760), .A1 (n_6_847), .A2 (slo___n23463));
NAND2_X1 slo__sro_c42890 (.ZN (slo__sro_n38759), .A1 (slo__sro_n38760), .A2 (slo__sro_n38761));
NAND2_X1 CLOCK_slo__sro_c59889 (.ZN (CLOCK_slo__sro_n54489), .A1 (n_6_2115), .A2 (n_6_1_203));
AOI21_X2 slo__sro_c43068 (.ZN (slo__sro_n38915), .A (slo__sro_n4313), .B1 (n_6_1264), .B2 (slo___n23274));
INV_X1 slo__c42916 (.ZN (slo__n38783), .A (n_6_1_883));
NAND2_X1 slo__sro_c43098 (.ZN (slo__sro_n38942), .A1 (n_6_1_204), .A2 (n_6_1690));
AND2_X2 slo__sro_c43069 (.ZN (slo__sro_n4312), .A1 (slo__sro_n38915), .A2 (slo__sro_n38916));
INV_X1 slo__sro_c43097 (.ZN (slo__sro_n38943), .A (slo__sro_n20081));
INV_X1 slo__c42986 (.ZN (slo__n38840), .A (n_6_1_165));
NAND2_X2 CLOCK_sgo__sro_c51365 (.ZN (CLOCK_sgo__sro_n47148), .A1 (CLOCK_sgo__sro_n47149), .A2 (CLOCK_sgo__sro_n47150));
NAND2_X1 slo__sro_c42947 (.ZN (slo__sro_n38808), .A1 (n_6_1_764), .A2 (n_6_668));
NAND2_X1 slo__sro_c42948 (.ZN (slo__sro_n38807), .A1 (slo__sro_n38808), .A2 (slo__sro_n12060));
AOI21_X2 slo__sro_c42949 (.ZN (n_6_1_759), .A (slo__sro_n38807), .B1 (n_6_700), .B2 (n_6_1_765));
INV_X2 slo__c43148 (.ZN (slo__n38973), .A (n_6_1_328));
INV_X32 CLOCK_slo__c67285 (.ZN (n_6_1_100), .A (CLOCK_slo__n60587));
AOI222_X2 CLOCK_slo__sro_c71859 (.ZN (CLOCK_slo__sro_n64581), .A1 (n_6_1893), .A2 (n_6_1_100)
    , .B1 (n_6_1861), .B2 (n_6_1_99), .C1 (opt_ipo_n24075), .C2 (n_6_1_98));
INV_X1 slo__c43601 (.ZN (slo__n39345), .A (CLOCK_slo__sro_n54789));
INV_X2 slo__c43277 (.ZN (slo__n39084), .A (n_6_1_929));
INV_X1 slo__c43341 (.ZN (slo__n39136), .A (slo__sro_n30017));
AND2_X1 CLOCK_slo__sro_c66505 (.ZN (CLOCK_slo__sro_n59951), .A1 (n_6_1582), .A2 (slo___n23244));
CLKBUF_X1 slo__L2_c2_c43529 (.Z (slo__n39284), .A (slo__n39285));
INV_X2 slo__c43691 (.ZN (slo__n39417), .A (slo__sro_n13471));
INV_X1 slo__c44054 (.ZN (slo__n39719), .A (slo__sro_n15534));
NAND2_X1 slo__sro_c44163 (.ZN (slo__sro_n39797), .A1 (n_6_1_150), .A2 (n_6_1_133));
AOI222_X2 slo__sro_c43893 (.ZN (slo__sro_n39597), .A1 (n_6_1446), .A2 (n_6_1_345)
    , .B1 (n_6_1414), .B2 (slo___n23229), .C1 (n_6_2238), .C2 (n_6_1_343));
AOI222_X2 slo__sro_c43854 (.ZN (slo__n39286), .A1 (n_6_1746), .A2 (n_6_1_169), .B1 (n_6_1778)
    , .B2 (CLOCK_sgo__n48020), .C1 (n_6_2095), .C2 (n_6_1_168));
NAND2_X1 CLOCK_slo__sro_c66704 (.ZN (CLOCK_slo__sro_n60127), .A1 (n_6_403), .A2 (n_6_1_904));
NAND2_X1 slo__sro_c44164 (.ZN (slo__sro_n39796), .A1 (n_6_1805), .A2 (n_6_1_134));
NAND2_X1 slo__sro_c44139 (.ZN (slo__sro_n39768), .A1 (n_0_59), .A2 (slo__sro_n39770));
INV_X1 opt_ipo_c28238 (.ZN (opt_ipo_n24861), .A (slo__sro_n29362));
INV_X1 slo__sro_c44137 (.ZN (slo__sro_n39770), .A (hfn_ipo_n33));
NAND2_X1 slo__sro_c44138 (.ZN (slo__sro_n39769), .A1 (slo__mro_n33299), .A2 (hfn_ipo_n33));
NOR2_X1 slo__sro_c44294 (.ZN (slo__sro_n39898), .A1 (slo__sro_n8415), .A2 (slo__sro_n39899));
NAND2_X1 slo__sro_c44414 (.ZN (slo__sro_n40009), .A1 (n_6_1413), .A2 (slo___n23229));
NAND2_X1 slo__sro_c44292 (.ZN (slo__sro_n39900), .A1 (n_6_82), .A2 (n_6_1_1079));
NAND2_X1 slo__sro_c44415 (.ZN (slo__sro_n40008), .A1 (slo__sro_n40009), .A2 (slo__sro_n40010));
INV_X1 CLOCK_sgo__sro_c51546 (.ZN (CLOCK_sgo__sro_n47298), .A (slo__sro_n29381));
AOI21_X2 slo__sro_c44416 (.ZN (slo__sro_n40007), .A (slo__sro_n40008), .B1 (n_6_1445), .B2 (n_6_1_345));
NAND2_X2 slo__sro_c46338 (.ZN (slo__sro_n41832), .A1 (n_6_251), .A2 (n_6_1_1010));
INV_X1 slo__c44354 (.ZN (slo__n39957), .A (slo__sro_n2346));
NAND2_X1 CLOCK_slo__sro_c53634 (.ZN (CLOCK_slo__sro_n49069), .A1 (slo___n16308), .A2 (n_6_1_868));
AND2_X2 slo__sro_c45537 (.ZN (n_6_1_684), .A1 (slo__sro_n41061), .A2 (slo__sro_n41060));
INV_X2 slo__c44107 (.ZN (slo__n39745), .A (n_6_1_129));
INV_X2 slo__c44505 (.ZN (slo__n40090), .A (n_6_1_96));
INV_X1 slo__sro_c45504 (.ZN (slo__sro_n41030), .A (slo__sro_n41031));
AND2_X1 slo__sro_c44729 (.ZN (slo__sro_n40292), .A1 (n_6_2383), .A2 (n_6_1_483));
AOI21_X1 slo__sro_c45503 (.ZN (slo__sro_n41031), .A (slo__sro_n7422), .B1 (n_6_996), .B2 (slo___n23218));
NAND2_X1 slo__sro_c46314 (.ZN (slo__sro_n41810), .A1 (n_6_2102), .A2 (n_6_1_168));
AOI21_X2 slo__sro_c45505 (.ZN (slo__sro_n41029), .A (slo__sro_n41030), .B1 (n_6_964), .B2 (slo___n23232));
NAND2_X1 slo__sro_c44578 (.ZN (slo__sro_n40150), .A1 (n_6_1_553), .A2 (n_6_2430));
NAND2_X1 slo__sro_c44579 (.ZN (slo__sro_n40149), .A1 (slo___n23457), .A2 (n_6_1068));
NAND2_X1 slo__sro_c44580 (.ZN (slo__sro_n40148), .A1 (slo__sro_n40149), .A2 (slo__sro_n40150));
INV_X1 CLOCK_slo__sro_c60593 (.ZN (CLOCK_slo__sro_n55087), .A (slo__sro_n22458));
AND2_X2 slo__sro_c45973 (.ZN (slo__sro_n41479), .A1 (n_6_1669), .A2 (slo___n23239));
NAND2_X1 slo__sro_c45535 (.ZN (slo__sro_n41061), .A1 (n_6_823), .A2 (n_6_1_695));
NAND2_X1 slo__sro_c45629 (.ZN (slo__sro_n41144), .A1 (n_6_2267), .A2 (n_6_1_378));
NAND2_X1 slo__sro_c44815 (.ZN (slo__sro_n40371), .A1 (n_6_2456), .A2 (n_6_1_588));
NAND2_X2 CLOCK_slo__mro_c70356 (.ZN (CLOCK_slo__mro_n63339), .A1 (n_6_1400), .A2 (n_6_1_380));
AND2_X1 CLOCK_slo__sro_c55215 (.ZN (CLOCK_slo__sro_n50484), .A1 (n_6_1460), .A2 (n_6_1_345));
BUF_X8 slo___L1_c47637 (.Z (slo___n43257), .A (n_6_1_415));
INV_X1 slo__sro_c45433 (.ZN (slo__sro_n40961), .A (n_6_1_798));
NOR2_X1 slo__sro_c45411 (.ZN (slo__sro_n40937), .A1 (slo__sro_n40939), .A2 (slo__sro_n40938));
AND2_X1 slo__sro_c45239 (.ZN (slo__sro_n40770), .A1 (n_6_2880), .A2 (CLOCK_sgo__n46945));
INV_X1 slo__sro_c44914 (.ZN (slo__sro_n40462), .A (slo__sro_n21603));
AOI222_X2 CLOCK_slo__sro_c71406 (.ZN (slo__sro_n39122), .A1 (n_6_1263), .A2 (slo___n23274)
    , .B1 (n_6_1231), .B2 (slo___n23359), .C1 (n_6_2340), .C2 (n_6_1_448));
NAND2_X2 slo__sro_c44916 (.ZN (slo__sro_n40460), .A1 (CLOCK_slo__mro_n63532), .A2 (slo__sro_n40462));
AOI21_X4 slo__sro_c44917 (.ZN (slo__sro_n40459), .A (slo__sro_n40460), .B1 (n_6_1299), .B2 (n_6_1_414));
CLKBUF_X1 CLOCK_slo___L1_c1_c72417 (.Z (n_6_2789), .A (CLOCK_slo___n65042));
AOI21_X2 slo__sro_c46317 (.ZN (slo__sro_n41807), .A (slo__sro_n41808), .B1 (n_6_1785), .B2 (CLOCK_sgo__n48020));
NAND2_X2 slo__sro_c46339 (.ZN (slo__sro_n41831), .A1 (slo__sro_n41832), .A2 (slo__sro_n41833));
INV_X2 opt_ipo_c28343 (.ZN (opt_ipo_n24966), .A (slo__sro_n9429));
AOI21_X2 CLOCK_slo__sro_c69412 (.ZN (slo__sro_n36308), .A (CLOCK_slo__sro_n62512)
    , .B1 (n_6_1378), .B2 (n_6_1_380));
NAND2_X2 slo__sro_c46316 (.ZN (slo__sro_n41808), .A1 (slo__sro_n41809), .A2 (slo__sro_n41810));
INV_X2 opt_ipo_c49477 (.ZN (opt_ipo_n45134), .A (n_6_1_444));
INV_X1 CLOCK_opt_ipo_c50150 (.ZN (CLOCK_opt_ipo_n45807), .A (n_6_1_419));
AOI21_X2 slo__sro_c46801 (.ZN (slo__sro_n42341), .A (CLOCK_slo__mro_n52173), .B1 (n_6_902), .B2 (slo___n23367));
NAND2_X1 CLOCK_sgo__sro_c51547 (.ZN (CLOCK_sgo__sro_n47297), .A1 (n_6_1486), .A2 (n_6_1_309));
NAND2_X1 CLOCK_sgo__sro_c51548 (.ZN (CLOCK_sgo__sro_n47296), .A1 (CLOCK_sgo__sro_n47297), .A2 (CLOCK_sgo__sro_n47298));
AOI21_X1 CLOCK_sgo__sro_c51549 (.ZN (slo__sro_n29380), .A (CLOCK_sgo__sro_n47296)
    , .B1 (n_6_1518), .B2 (slo___n23247));
NAND2_X1 CLOCK_sgo__sro_c51559 (.ZN (CLOCK_sgo__sro_n47307), .A1 (opt_ipo_n24173), .A2 (n_6_1_868));
INV_X1 CLOCK_slo__sro_c69830 (.ZN (CLOCK_slo__sro_n62895), .A (slo__sro_n40770));
AOI21_X1 CLOCK_slo__sro_c65776 (.ZN (CLOCK_slo__sro_n59280), .A (CLOCK_slo__sro_n59281)
    , .B1 (n_6_206), .B2 (n_6_1_1009));
INV_X4 CLOCK_opt_ipo_c50122 (.ZN (CLOCK_opt_ipo_n45779), .A (slo__sro_n32470));
INV_X1 opt_ipo_c48278 (.ZN (opt_ipo_n43935), .A (slo__sro_n28333));
BUF_X2 spt__c74549 (.Z (n_6_1_305), .A (spt__n66340));
BUF_X8 CLOCK_sgo__L2_c2_c51054 (.Z (CLOCK_sgo__n46814), .A (CLOCK_sgo__n46815));
INV_X1 CLOCK_opt_ipo_c50168 (.ZN (CLOCK_opt_ipo_n45825), .A (n_6_1_523));
INV_X4 opt_ipo_c28383 (.ZN (opt_ipo_n25006), .A (opt_ipo_n25007));
BUF_X4 opt_ipo_c28384 (.Z (opt_ipo_n25007), .A (n_6_1_1006));
NAND2_X1 CLOCK_sgo__sro_c51664 (.ZN (CLOCK_sgo__sro_n47394), .A1 (CLOCK_sgo__sro_n47395), .A2 (slo__sro_n21678));
AOI21_X4 CLOCK_sgo__sro_c51665 (.ZN (slo__sro_n21676), .A (CLOCK_sgo__sro_n47394)
    , .B1 (n_6_706), .B2 (n_6_1_729));
BUF_X4 CLOCK_sgo__L1_c1_c51055 (.Z (CLOCK_sgo__n46815), .A (drc_ipoPP_2PP_0));
INV_X4 opt_ipo_c49487 (.ZN (opt_ipo_n45144), .A (opt_ipo_n45145));
AOI21_X4 CLOCK_sgo__sro_c51438 (.ZN (slo__sro_n19627), .A (CLOCK_sgo__sro_n47210)
    , .B1 (n_6_1528), .B2 (slo___n23247));
NAND2_X1 CLOCK_sgo__sro_c51592 (.ZN (CLOCK_sgo__sro_n47338), .A1 (n_6_614), .A2 (n_6_1_800));
BUF_X2 opt_ipo_c49488 (.Z (opt_ipo_n45145), .A (n_6_1_516));
NAND2_X1 CLOCK_sgo__sro_c51593 (.ZN (CLOCK_sgo__sro_n47337), .A1 (CLOCK_sgo__sro_n47338), .A2 (CLOCK_sgo__sro_n47339));
BUF_X1 slo___L1_c47627 (.Z (slo___n43247), .A (n_6_1_100));
NAND2_X1 CLOCK_sgo__sro_c51424 (.ZN (CLOCK_sgo__sro_n47198), .A1 (CLOCK_sgo__sro_n47199), .A2 (CLOCK_sgo__sro_n47200));
AOI21_X2 CLOCK_sgo__sro_c51425 (.ZN (CLOCK_sgo__sro_n47197), .A (CLOCK_sgo__sro_n47198)
    , .B1 (n_6_324), .B2 (n_6_1_939));
INV_X1 CLOCK_sgo__sro_c51785 (.ZN (CLOCK_sgo__sro_n47503), .A (slo__sro_n35250));
NAND2_X1 CLOCK_sgo__sro_c51786 (.ZN (CLOCK_sgo__sro_n47502), .A1 (n_6_646), .A2 (n_6_1_764));
INV_X1 CLOCK_sgo__sro_c51716 (.ZN (CLOCK_sgo__sro_n47442), .A (slo__sro_n5946));
NAND2_X1 CLOCK_sgo__sro_c51717 (.ZN (CLOCK_sgo__sro_n47441), .A1 (n_6_1_379), .A2 (n_6_1349));
INV_X1 CLOCK_sgo__sro_c51435 (.ZN (CLOCK_sgo__sro_n47212), .A (slo__sro_n19628));
BUF_X8 CLOCK_sgo__L1_c1_c51064 (.Z (drc_ipo_n26621), .A (CLOCK_sgo__n46841));
NAND2_X2 CLOCK_sgo__sro_c51436 (.ZN (CLOCK_sgo__sro_n47211), .A1 (n_6_1496), .A2 (n_6_1_309));
INV_X4 CLOCK_opt_ipo_c50146 (.ZN (CLOCK_opt_ipo_n45803), .A (slo__sro_n6673));
NAND2_X1 CLOCK_sgo__sro_c51718 (.ZN (CLOCK_sgo__sro_n47440), .A1 (CLOCK_sgo__sro_n47441), .A2 (CLOCK_sgo__sro_n47442));
AOI21_X2 CLOCK_sgo__sro_c51719 (.ZN (slo__sro_n5945), .A (CLOCK_sgo__sro_n47440), .B1 (n_6_1381), .B2 (n_6_1_380));
AOI21_X1 CLOCK_sgo__sro_c51788 (.ZN (slo__sro_n35249), .A (CLOCK_sgo__sro_n47501)
    , .B1 (n_6_678), .B2 (n_6_1_765));
INV_X1 CLOCK_sgo__sro_c51836 (.ZN (CLOCK_sgo__sro_n47540), .A (n_6_1_134));
NAND2_X1 CLOCK_sgo__sro_c51837 (.ZN (CLOCK_sgo__sro_n47539), .A1 (n_6_2054), .A2 (n_6_1_133));
AOI21_X1 CLOCK_sgo__sro_c51864 (.ZN (n_6_1_911), .A (CLOCK_sgo__sro_n47560), .B1 (n_6_325), .B2 (n_6_1_939));
OAI21_X1 CLOCK_sgo__sro_c51838 (.ZN (CLOCK_sgo__sro_n47538), .A (CLOCK_sgo__sro_n47539)
    , .B1 (CLOCK_sgo__sro_n47541), .B2 (CLOCK_sgo__sro_n47540));
AOI21_X1 CLOCK_sgo__sro_c51839 (.ZN (n_6_1_109), .A (CLOCK_sgo__sro_n47538), .B1 (n_6_1832), .B2 (n_6_1_135));
INV_X1 CLOCK_sgo__sro_c51861 (.ZN (CLOCK_sgo__sro_n47562), .A (slo__sro_n11080));
NAND2_X1 CLOCK_sgo__sro_c51862 (.ZN (CLOCK_sgo__sro_n47561), .A1 (n_6_357), .A2 (n_6_1_940));
INV_X4 CLOCK_opt_ipo_c50216 (.ZN (CLOCK_opt_ipo_n45873), .A (slo__sro_n14522));
NAND2_X2 CLOCK_sgo__sro_c51911 (.ZN (CLOCK_sgo__sro_n47603), .A1 (n_6_1814), .A2 (n_6_1_134));
NAND2_X1 CLOCK_sgo__sro_c51912 (.ZN (CLOCK_sgo__sro_n47602), .A1 (CLOCK_sgo__sro_n47603), .A2 (CLOCK_sgo__sro_n47604));
AOI21_X1 CLOCK_sgo__sro_c51913 (.ZN (n_6_1_123), .A (CLOCK_sgo__sro_n47602), .B1 (n_6_1846), .B2 (n_6_1_135));
INV_X1 CLOCK_sgo__sro_c51933 (.ZN (CLOCK_sgo__sro_n47623), .A (slo__sro_n28681));
NAND2_X1 CLOCK_sgo__sro_c51934 (.ZN (CLOCK_sgo__sro_n47622), .A1 (n_6_1618), .A2 (slo___n23215));
NAND2_X1 CLOCK_sgo__sro_c51935 (.ZN (CLOCK_sgo__sro_n47621), .A1 (CLOCK_sgo__sro_n47622), .A2 (CLOCK_sgo__sro_n47623));
AOI21_X2 CLOCK_sgo__sro_c51936 (.ZN (n_6_1_224), .A (CLOCK_sgo__sro_n47621), .B1 (n_6_1650), .B2 (drc_ipo_n26601));
AOI21_X2 CLOCK_sgo__sro_c51985 (.ZN (slo__sro_n10712), .A (CLOCK_sgo__sro_n47663)
    , .B1 (n_6_1640), .B2 (drc_ipo_n26601));
INV_X2 CLOCK_opt_ipo_c50236 (.ZN (CLOCK_opt_ipo_n45893), .A (CLOCK_opt_ipo_n45894));
BUF_X2 CLOCK_opt_ipo_c50237 (.Z (CLOCK_opt_ipo_n45894), .A (CLOCK_slo__sro_n59549));
NAND2_X1 CLOCK_slo__sro_c68485 (.ZN (CLOCK_slo__sro_n61698), .A1 (n_6_2887), .A2 (slo__n13799));
INV_X1 CLOCK_sgo__sro_c52006 (.ZN (CLOCK_sgo__sro_n47682), .A (CLOCK_sgo__sro_n47683));
AOI221_X2 CLOCK_sgo__sro_c52007 (.ZN (n_6_1_243), .A (CLOCK_sgo__sro_n47682), .B1 (n_6_1538)
    , .B2 (n_6_1_274), .C1 (n_6_1570), .C2 (slo___n23244));
AOI221_X2 CLOCK_sgo__sro_c52038 (.ZN (n_6_1_212), .A (CLOCK_sgo__sro_n47701), .B1 (n_6_1606)
    , .B2 (slo___n23215), .C1 (n_6_1638), .C2 (drc_ipo_n26601));
INV_X1 CLOCK_opt_ipo_c50079 (.ZN (CLOCK_opt_ipo_n45736), .A (slo__sro_n13037));
INV_X4 opt_ipo_c28493 (.ZN (opt_ipo_n25116), .A (slo__sro_n21753));
INV_X4 CLOCK_opt_ipo_c50249 (.ZN (CLOCK_opt_ipo_n45906), .A (n_6_1_384));
INV_X1 opt_ipo_c28497 (.ZN (opt_ipo_n25120), .A (n_6_1_985));
NAND2_X2 CLOCK_sgo__sro_c51310 (.ZN (CLOCK_sgo__sro_n47110), .A1 (n_6_1752), .A2 (n_6_1_169));
NAND2_X1 CLOCK_slo__sro_c68050 (.ZN (CLOCK_slo__sro_n61283), .A1 (CLOCK_slo__sro_n61284), .A2 (slo__sro_n3862));
NAND2_X1 CLOCK_sgo__sro_c52080 (.ZN (CLOCK_sgo__sro_n47733), .A1 (n_6_1_309), .A2 (n_6_1477));
INV_X2 CLOCK_opt_ipo_c50261 (.ZN (CLOCK_opt_ipo_n45918), .A (n_6_1_452));
AOI21_X2 CLOCK_slo__sro_c68051 (.ZN (slo__sro_n3860), .A (CLOCK_slo__sro_n61283), .B1 (n_6_1452), .B2 (n_6_1_345));
BUF_X2 CLOCK_sgo__c51165 (.Z (n_6_1_973), .A (CLOCK_sgo__n46942));
INV_X2 CLOCK_slo__c53090 (.ZN (slo__sro_n34940), .A (CLOCK_slo__n48588));
NAND2_X1 CLOCK_slo__sro_c68587 (.ZN (CLOCK_slo__sro_n61785), .A1 (n_6_1_134), .A2 (n_6_1797));
INV_X1 CLOCK_sgo__sro_c52161 (.ZN (CLOCK_sgo__sro_n47801), .A (slo__sro_n5027));
INV_X2 opt_ipo_c48448 (.ZN (opt_ipo_n44105), .A (n_6_1_862));
INV_X1 CLOCK_slo__sro_c68125 (.ZN (CLOCK_slo__sro_n61348), .A (CLOCK_slo__sro_n61349));
NAND2_X1 CLOCK_sgo__sro_c52114 (.ZN (CLOCK_sgo__sro_n47761), .A1 (n_6_1_379), .A2 (n_6_1351));
NAND2_X1 CLOCK_sgo__sro_c52115 (.ZN (CLOCK_sgo__sro_n47760), .A1 (CLOCK_sgo__sro_n47761), .A2 (CLOCK_sgo__sro_n47762));
AOI21_X2 CLOCK_sgo__sro_c52116 (.ZN (slo__sro_n20146), .A (CLOCK_sgo__sro_n47760)
    , .B1 (n_6_1383), .B2 (n_6_1_380));
INV_X1 opt_ipo_c48459 (.ZN (opt_ipo_n44116), .A (CLOCK_slo__sro_n60679));
AOI21_X4 CLOCK_sgo__sro_c52164 (.ZN (CLOCK_sgo__sro_n47798), .A (CLOCK_sgo__sro_n47799)
    , .B1 (n_6_1403), .B2 (n_6_1_380));
AOI221_X2 CLOCK_slo__sro_c52820 (.ZN (slo__sro_n35163), .A (CLOCK_slo__sro_n48338)
    , .B1 (n_6_645), .B2 (n_6_1_764), .C1 (n_6_677), .C2 (n_6_1_765));
NAND2_X4 CLOCK_slo__mro_c53131 (.ZN (slo__sro_n8604), .A1 (n_6_98), .A2 (n_6_1_1080));
INV_X1 CLOCK_sgo__sro_c52191 (.ZN (CLOCK_sgo__sro_n47825), .A (slo__sro_n15657));
NAND2_X1 CLOCK_sgo__sro_c52192 (.ZN (CLOCK_sgo__sro_n47824), .A1 (n_6_1497), .A2 (n_6_1_309));
NAND2_X2 CLOCK_sgo__sro_c52193 (.ZN (CLOCK_sgo__sro_n47823), .A1 (CLOCK_sgo__sro_n47824), .A2 (CLOCK_sgo__sro_n47825));
AOI21_X4 CLOCK_sgo__sro_c52194 (.ZN (CLOCK_sgo__sro_n47822), .A (CLOCK_sgo__sro_n47823)
    , .B1 (n_6_1529), .B2 (slo___n23247));
NAND2_X1 CLOCK_sgo__sro_c52204 (.ZN (CLOCK_sgo__sro_n47837), .A1 (n_6_1275), .A2 (slo___n23274));
AOI21_X1 CLOCK_sgo__sro_c52205 (.ZN (CLOCK_sgo__sro_n47836), .A (slo__sro_n11889)
    , .B1 (n_6_1243), .B2 (slo___n23359));
AND2_X2 CLOCK_sgo__sro_c52206 (.ZN (CLOCK_sgo__sro_n47835), .A1 (CLOCK_sgo__sro_n47837), .A2 (CLOCK_sgo__sro_n47836));
INV_X4 CLOCK_opt_ipo_c50312 (.ZN (CLOCK_opt_ipo_n45969), .A (slo__sro_n6160));
AOI21_X1 CLOCK_sgo__sro_c52216 (.ZN (CLOCK_sgo__sro_n47846), .A (slo__sro_n2969), .B1 (n_6_1434), .B2 (slo___n23229));
INV_X1 CLOCK_sgo__sro_c52503 (.ZN (CLOCK_sgo__sro_n48087), .A (slo__sro_n11858));
INV_X4 CLOCK_opt_ipo_c50321 (.ZN (CLOCK_opt_ipo_n45978), .A (n_6_1_354));
INV_X2 opt_ipo_c49709 (.ZN (opt_ipo_n45366), .A (n_6_1_616));
NAND2_X2 CLOCK_sgo__sro_c52505 (.ZN (CLOCK_sgo__sro_n48085), .A1 (CLOCK_sgo__sro_n48086), .A2 (CLOCK_sgo__sro_n48087));
AOI21_X4 CLOCK_sgo__sro_c52506 (.ZN (n_6_1_943), .A (CLOCK_sgo__sro_n48085), .B1 (n_6_258), .B2 (n_6_1_974));
NAND2_X1 CLOCK_sgo__sro_c52625 (.ZN (CLOCK_sgo__sro_n48189), .A1 (CLOCK_sgo__sro_n48190), .A2 (slo__sro_n32140));
BUF_X8 CLOCK_sgo__L2_c2_c51218 (.Z (n_6_17), .A (CLOCK_sgo__n47004));
AOI21_X1 CLOCK_slo__sro_c68795 (.ZN (slo__sro_n9268), .A (CLOCK_slo__sro_n61961), .B1 (n_6_1168), .B2 (slo___n23364));
CLKBUF_X3 CLOCK_sgo__L1_c3_c51220 (.Z (CLOCK_sgo__n47002), .A (CLOCK_sgo__n47005));
AOI21_X2 CLOCK_sgo__sro_c52626 (.ZN (slo__sro_n32138), .A (CLOCK_sgo__sro_n48189)
    , .B1 (n_6_322), .B2 (n_6_1_939));
NAND2_X1 CLOCK_slo__sro_c53265 (.ZN (CLOCK_slo__sro_n48740), .A1 (CLOCK_slo__sro_n48741), .A2 (CLOCK_slo__sro_n48742));
AOI21_X2 CLOCK_slo__sro_c53266 (.ZN (n_6_1_213), .A (CLOCK_slo__sro_n48740), .B1 (n_6_1639), .B2 (drc_ipo_n26601));
NAND2_X1 CLOCK_slo__sro_c53348 (.ZN (CLOCK_slo__sro_n48814), .A1 (n_6_1358), .A2 (n_6_1_379));
INV_X1 CLOCK_opt_ipo_c50348 (.ZN (CLOCK_opt_ipo_n46005), .A (n_6_1_567));
INV_X1 CLOCK_slo__sro_c53416 (.ZN (CLOCK_slo__sro_n48876), .A (slo___n8747));
NAND2_X2 CLOCK_slo__mro_c69068 (.ZN (CLOCK_slo__mro_n62209), .A1 (n_6_1701), .A2 (slo___n23407));
NAND2_X1 CLOCK_slo__sro_c68982 (.ZN (CLOCK_slo__sro_n62130), .A1 (n_6_237), .A2 (n_6_1_1010));
NAND2_X1 CLOCK_slo__sro_c68983 (.ZN (CLOCK_slo__sro_n62129), .A1 (CLOCK_slo__sro_n62130), .A2 (CLOCK_slo__sro_n62131));
NOR2_X2 CLOCK_slo__sro_c69204 (.ZN (n_6_1_371), .A1 (CLOCK_sgo__sro_n47134), .A2 (CLOCK_slo__sro_n62332));
INV_X1 CLOCK_slo__sro_c53417 (.ZN (CLOCK_slo__sro_n48875), .A (n_6_1_868));
NAND2_X1 CLOCK_slo__sro_c53349 (.ZN (CLOCK_slo__sro_n48813), .A1 (CLOCK_slo__sro_n48814), .A2 (CLOCK_slo__sro_n48815));
NAND2_X1 CLOCK_slo__sro_c53318 (.ZN (CLOCK_slo__sro_n48786), .A1 (slo___n15724), .A2 (n_6_1_308));
INV_X1 CLOCK_slo__sro_c53319 (.ZN (CLOCK_slo__sro_n48785), .A (CLOCK_slo__sro_n48786));
NAND2_X2 CLOCK_slo__mro_c70808 (.ZN (slo__sro_n7774), .A1 (n_6_228), .A2 (n_6_1_1010));
INV_X2 CLOCK_opt_ipo_c50372 (.ZN (CLOCK_opt_ipo_n46029), .A (slo__sro_n37192));
NOR2_X1 CLOCK_slo__sro_c53418 (.ZN (CLOCK_slo__sro_n48874), .A1 (CLOCK_slo__sro_n48876), .A2 (CLOCK_slo__sro_n48875));
AOI221_X2 CLOCK_slo__sro_c53419 (.ZN (slo__sro_n8731), .A (CLOCK_slo__sro_n48874)
    , .B1 (n_6_457), .B2 (n_6_1_869), .C1 (n_6_489), .C2 (n_6_1_870));
AOI21_X2 CLOCK_slo__sro_c53511 (.ZN (slo__sro_n13461), .A (CLOCK_slo__sro_n48958)
    , .B1 (n_6_1483), .B2 (n_6_1_309));
INV_X2 CLOCK_opt_ipo_c50381 (.ZN (CLOCK_opt_ipo_n46038), .A (slo__sro_n8731));
NAND2_X1 CLOCK_slo__sro_c53532 (.ZN (CLOCK_slo__sro_n48976), .A1 (CLOCK_slo__sro_n48977), .A2 (CLOCK_slo__sro_n48978));
AOI21_X2 CLOCK_slo__sro_c53533 (.ZN (n_6_1_112), .A (CLOCK_slo__sro_n48976), .B1 (n_6_1835), .B2 (n_6_1_135));
BUF_X4 CLOCK_sgo__L2_c2_c51259 (.Z (n_6_23), .A (CLOCK_sgo__n47049));
BUF_X2 CLOCK_sgo__L1_c1_c51260 (.Z (CLOCK_sgo__n47049), .A (CLOCK_sgo__n47051));
BUF_X8 CLOCK_sgo__L1_c1_c51261 (.Z (drc_ipo_n26575), .A (CLOCK_sgo__n47054));
NAND2_X1 CLOCK_slo__sro_c53582 (.ZN (CLOCK_slo__sro_n49024), .A1 (n_6_1179), .A2 (slo___n23364));
NAND2_X1 CLOCK_slo__sro_c53583 (.ZN (CLOCK_slo__sro_n49023), .A1 (CLOCK_slo__sro_n49025), .A2 (CLOCK_slo__sro_n49024));
AOI21_X2 CLOCK_slo__sro_c53584 (.ZN (CLOCK_slo__sro_n49022), .A (CLOCK_slo__sro_n49023)
    , .B1 (n_6_1211), .B2 (slo___n23466));
INV_X2 CLOCK_slo__c53616 (.ZN (n_6_1_734), .A (CLOCK_slo__n49050));
NAND2_X1 CLOCK_slo__sro_c69712 (.ZN (CLOCK_slo__sro_n62785), .A1 (n_6_846), .A2 (slo___n23463));
AOI221_X2 CLOCK_slo__sro_c53655 (.ZN (slo__sro_n17693), .A (CLOCK_slo__sro_n49084)
    , .B1 (n_6_1255), .B2 (slo___n23274), .C1 (n_6_1223), .C2 (slo___n23359));
INV_X1 CLOCK_slo__sro_c53695 (.ZN (CLOCK_slo__sro_n49120), .A (CLOCK_slo__sro_n49121));
AOI221_X2 CLOCK_slo__sro_c53696 (.ZN (n_6_1_601), .A (CLOCK_slo__sro_n49120), .B1 (n_6_906)
    , .B2 (slo___n23367), .C1 (n_6_938), .C2 (n_6_1_625));
INV_X32 CLOCK_slo__c53719 (.ZN (n_6_1_414), .A (CLOCK_slo__n49141));
NAND2_X1 CLOCK_slo__sro_c53772 (.ZN (CLOCK_slo__sro_n49191), .A1 (n_6_1_798), .A2 (n_6_2649));
NAND2_X1 CLOCK_slo__sro_c53773 (.ZN (CLOCK_slo__sro_n49190), .A1 (n_6_622), .A2 (n_6_1_800));
AOI21_X1 CLOCK_slo__sro_c68173 (.ZN (CLOCK_slo__sro_n61395), .A (slo__sro_n5017), .B1 (n_6_1301), .B2 (n_6_1_414));
INV_X4 opt_ipo_c49823 (.ZN (CLOCK_spw__n65836), .A (n_6_1_1081));
INV_X1 CLOCK_slo__sro_c53801 (.ZN (CLOCK_slo__sro_n49218), .A (n_6_2707));
INV_X1 CLOCK_slo__sro_c53802 (.ZN (CLOCK_slo__sro_n49217), .A (n_6_1_868));
NOR2_X1 CLOCK_slo__sro_c53803 (.ZN (CLOCK_slo__sro_n49216), .A1 (CLOCK_slo__sro_n49218), .A2 (CLOCK_slo__sro_n49217));
AOI222_X1 CLOCK_slo__sro_c64754 (.ZN (n_6_1_976), .A1 (n_6_224), .A2 (n_6_1_1010)
    , .B1 (n_6_192), .B2 (n_6_1_1009), .C1 (n_6_2821), .C2 (CLOCK_sgo__n46950));
CLKBUF_X2 spt__c74604 (.Z (CLOCK_sgo__sro_n47592), .A (spt__n66402));
NAND2_X1 CLOCK_slo__sro_c53956 (.ZN (CLOCK_slo__sro_n49349), .A1 (slo___n23229), .A2 (n_6_1427));
NAND2_X1 CLOCK_slo__sro_c53957 (.ZN (CLOCK_slo__sro_n49348), .A1 (CLOCK_slo__sro_n49349), .A2 (CLOCK_slo__sro_n49350));
AOI21_X2 CLOCK_slo__sro_c53958 (.ZN (n_6_1_330), .A (CLOCK_slo__sro_n49348), .B1 (n_6_1459), .B2 (n_6_1_345));
INV_X2 CLOCK_slo__sro_c53999 (.ZN (CLOCK_slo__sro_n49386), .A (n_6_801));
INV_X1 CLOCK_slo__sro_c54000 (.ZN (CLOCK_slo__sro_n49385), .A (n_6_1_695));
NAND2_X1 CLOCK_slo__sro_c54001 (.ZN (CLOCK_slo__sro_n49384), .A1 (n_6_2543), .A2 (n_6_1_693));
OAI21_X2 CLOCK_slo__sro_c54002 (.ZN (CLOCK_slo__sro_n49383), .A (CLOCK_slo__sro_n49384)
    , .B1 (CLOCK_slo__sro_n49386), .B2 (CLOCK_slo__sro_n49385));
AOI21_X2 CLOCK_slo__sro_c54003 (.ZN (CLOCK_slo__sro_n49382), .A (CLOCK_slo__sro_n49383)
    , .B1 (n_6_769), .B2 (n_6_1_694));
NAND2_X1 CLOCK_slo__sro_c54023 (.ZN (CLOCK_slo__sro_n49403), .A1 (n_6_1288), .A2 (n_6_1_414));
NAND2_X1 CLOCK_slo__sro_c54024 (.ZN (CLOCK_slo__sro_n49402), .A1 (CLOCK_slo__sro_n49403), .A2 (slo__sro_n9561));
INV_X2 CLOCK_opt_ipo_c50461 (.ZN (CLOCK_opt_ipo_n46124), .A (n_6_1_875));
NAND2_X1 CLOCK_slo__sro_c54052 (.ZN (CLOCK_slo__sro_n49428), .A1 (n_6_1_870), .A2 (n_6_496));
NAND2_X1 CLOCK_slo__sro_c56121 (.ZN (CLOCK_slo__sro_n51308), .A1 (n_6_142), .A2 (n_6_1_1044));
AOI21_X2 CLOCK_slo__sro_c54054 (.ZN (CLOCK_slo__sro_n49426), .A (CLOCK_slo__sro_n49427)
    , .B1 (n_6_464), .B2 (n_6_1_869));
INV_X1 CLOCK_opt_ipo_c50470 (.ZN (CLOCK_opt_ipo_n46133), .A (CLOCK_slo__sro_n55447));
AOI21_X4 CLOCK_slo__sro_c54230 (.ZN (CLOCK_slo__sro_n49602), .A (CLOCK_slo__sro_n49603)
    , .B1 (n_6_504), .B2 (n_6_1_870));
INV_X4 CLOCK_opt_ipo_c50474 (.ZN (CLOCK_opt_ipo_n46137), .A (slo__sro_n35270));
NAND2_X1 CLOCK_slo__sro_c54292 (.ZN (CLOCK_slo__sro_n49663), .A1 (n_6_1_379), .A2 (n_6_1352));
NAND2_X1 CLOCK_slo__sro_c54293 (.ZN (CLOCK_slo__sro_n49662), .A1 (CLOCK_slo__sro_n49663), .A2 (CLOCK_slo__sro_n49664));
AOI21_X2 CLOCK_slo__sro_c54294 (.ZN (n_6_1_354), .A (CLOCK_slo__sro_n49662), .B1 (n_6_1384), .B2 (n_6_1_380));
INV_X4 CLOCK_opt_ipo_c50483 (.ZN (CLOCK_opt_ipo_n46146), .A (slo__sro_n2106));
INV_X1 opt_ipo_c49899 (.ZN (opt_ipo_n45556), .A (n_6_537));
NAND2_X2 CLOCK_slo__sro_c54350 (.ZN (CLOCK_slo__sro_n49712), .A1 (CLOCK_slo__sro_n49713), .A2 (CLOCK_slo__sro_n49714));
AOI21_X4 CLOCK_slo__sro_c54351 (.ZN (slo__sro_n11383), .A (CLOCK_slo__sro_n49712)
    , .B1 (n_6_1161), .B2 (slo___n23364));
NAND2_X1 CLOCK_slo__sro_c54367 (.ZN (CLOCK_slo__sro_n49727), .A1 (slo___n23215), .A2 (n_6_1630));
INV_X2 opt_ipo_c49908 (.ZN (opt_ipo_n45565), .A (n_6_1_966));
AOI21_X2 CLOCK_slo__sro_c54369 (.ZN (n_6_1_236), .A (CLOCK_slo__sro_n49726), .B1 (n_6_1662), .B2 (drc_ipo_n26601));
NAND2_X1 CLOCK_slo__sro_c54403 (.ZN (CLOCK_slo__sro_n49760), .A1 (n_6_1_379), .A2 (n_6_1350));
NAND2_X2 CLOCK_slo__sro_c54404 (.ZN (CLOCK_slo__sro_n49759), .A1 (CLOCK_slo__sro_n49760), .A2 (CLOCK_slo__sro_n49761));
AOI21_X2 CLOCK_slo__sro_c68488 (.ZN (slo__sro_n34136), .A (CLOCK_slo__sro_n61696)
    , .B1 (n_6_100), .B2 (n_6_1_1080));
AOI21_X2 CLOCK_slo__sro_c54405 (.ZN (CLOCK_slo__sro_n49758), .A (CLOCK_slo__sro_n49759)
    , .B1 (n_6_1382), .B2 (n_6_1_380));
INV_X4 opt_ipo_c28771 (.ZN (opt_ipo_n25394), .A (n_6_1_601));
NAND2_X1 CLOCK_slo__sro_c54418 (.ZN (CLOCK_slo__sro_n49773), .A1 (CLOCK_slo__sro_n49774), .A2 (CLOCK_slo__sro_n49775));
AOI221_X2 CLOCK_slo__sro_c68126 (.ZN (CLOCK_slo__sro_n61347), .A (CLOCK_slo__sro_n61348)
    , .B1 (n_6_129), .B2 (n_6_1_1044), .C1 (n_6_161), .C2 (n_6_1_1045));
AOI21_X2 CLOCK_slo__sro_c54419 (.ZN (CLOCK_slo__sro_n49772), .A (CLOCK_slo__sro_n49773)
    , .B1 (n_6_1192), .B2 (slo___n23466));
NOR2_X2 CLOCK_slo__sro_c54514 (.ZN (n_6_1_1072), .A1 (slo__sro_n4814), .A2 (CLOCK_slo__sro_n49853));
NAND2_X1 CLOCK_slo__sro_c54528 (.ZN (CLOCK_slo__sro_n49864), .A1 (n_6_980), .A2 (slo___n23232));
INV_X2 CLOCK_opt_ipo_c50526 (.ZN (CLOCK_opt_ipo_n46189), .A (sgo__sro_n1559));
AOI21_X2 CLOCK_slo__sro_c54530 (.ZN (slo__sro_n6088), .A (CLOCK_slo__sro_n49863), .B1 (n_6_1012), .B2 (slo___n23218));
NAND2_X1 CLOCK_slo__sro_c54583 (.ZN (CLOCK_slo__sro_n49912), .A1 (n_6_1629), .A2 (slo___n23215));
NAND2_X1 CLOCK_slo__sro_c54584 (.ZN (CLOCK_slo__sro_n49911), .A1 (CLOCK_slo__sro_n49912), .A2 (CLOCK_slo__sro_n49913));
AOI21_X2 CLOCK_slo__sro_c54585 (.ZN (n_6_1_235), .A (CLOCK_slo__sro_n49911), .B1 (n_6_1661), .B2 (drc_ipo_n26601));
INV_X1 CLOCK_slo__sro_c54616 (.ZN (CLOCK_slo__sro_n49938), .A (n_6_1_98));
NOR2_X1 CLOCK_slo__sro_c54617 (.ZN (CLOCK_slo__sro_n49937), .A1 (CLOCK_slo__sro_n49939), .A2 (CLOCK_slo__sro_n49938));
INV_X1 opt_ipo_c48737 (.ZN (opt_ipo_n44394), .A (CLOCK_slo__sro_n58313));
NAND2_X1 CLOCK_slo__sro_c69832 (.ZN (CLOCK_slo__sro_n62893), .A1 (CLOCK_slo__sro_n62894), .A2 (CLOCK_slo__sro_n62895));
NAND2_X1 CLOCK_slo__sro_c54644 (.ZN (CLOCK_slo__sro_n49962), .A1 (n_6_1556), .A2 (n_6_1_274));
NAND2_X1 CLOCK_slo__sro_c54645 (.ZN (CLOCK_slo__sro_n49961), .A1 (CLOCK_slo__sro_n49962), .A2 (slo__sro_n6899));
AOI21_X2 CLOCK_slo__sro_c54646 (.ZN (slo__sro_n6897), .A (CLOCK_slo__sro_n49961), .B1 (n_6_1588), .B2 (slo___n23244));
INV_X1 CLOCK_slo__sro_c54758 (.ZN (CLOCK_slo__sro_n50071), .A (slo__sro_n10905));
NAND2_X1 CLOCK_slo__sro_c54759 (.ZN (CLOCK_slo__sro_n50070), .A1 (n_6_268), .A2 (n_6_1_974));
NAND2_X1 CLOCK_slo__sro_c54760 (.ZN (CLOCK_slo__sro_n50069), .A1 (CLOCK_slo__sro_n50070), .A2 (CLOCK_slo__sro_n50071));
AOI21_X2 CLOCK_slo__sro_c54761 (.ZN (CLOCK_slo__sro_n50068), .A (CLOCK_slo__sro_n50069)
    , .B1 (n_6_300), .B2 (n_6_1_975));
AOI21_X1 CLOCK_slo__sro_c54787 (.ZN (CLOCK_slo__sro_n50097), .A (slo__sro_n5075), .B1 (n_6_1418), .B2 (slo___n23229));
AND2_X2 CLOCK_slo__sro_c54788 (.ZN (CLOCK_slo__sro_n50096), .A1 (CLOCK_slo__sro_n50097), .A2 (CLOCK_slo__sro_n50098));
INV_X1 CLOCK_slo__sro_c54821 (.ZN (CLOCK_slo__sro_n50130), .A (CLOCK_slo__sro_n50131));
AOI221_X1 CLOCK_slo__sro_c54822 (.ZN (n_6_1_567), .A (CLOCK_slo__sro_n50130), .B1 (n_6_971)
    , .B2 (slo___n23232), .C1 (n_6_1003), .C2 (slo___n23218));
NAND2_X1 CLOCK_slo__sro_c54833 (.ZN (CLOCK_slo__sro_n50140), .A1 (n_6_1365), .A2 (n_6_1_379));
NAND2_X1 CLOCK_slo__sro_c54834 (.ZN (CLOCK_slo__sro_n50139), .A1 (CLOCK_slo__sro_n50140), .A2 (CLOCK_slo__sro_n50141));
AOI21_X2 CLOCK_slo__sro_c54835 (.ZN (CLOCK_slo__sro_n50138), .A (CLOCK_slo__sro_n50139)
    , .B1 (n_6_1397), .B2 (n_6_1_380));
NAND2_X2 CLOCK_slo__sro_c54884 (.ZN (CLOCK_slo__sro_n50187), .A1 (n_6_867), .A2 (n_6_1_660));
NAND2_X2 CLOCK_slo__sro_c54885 (.ZN (CLOCK_slo__sro_n50186), .A1 (CLOCK_slo__sro_n50187), .A2 (CLOCK_slo__sro_n50188));
AOI21_X2 CLOCK_slo__sro_c54886 (.ZN (n_6_1_629), .A (CLOCK_slo__sro_n50186), .B1 (n_6_835), .B2 (slo___n23463));
NAND2_X1 CLOCK_slo__sro_c54926 (.ZN (CLOCK_slo__sro_n50226), .A1 (n_6_1488), .A2 (n_6_1_309));
NAND2_X1 CLOCK_slo__sro_c54927 (.ZN (CLOCK_slo__sro_n50225), .A1 (CLOCK_slo__sro_n50226), .A2 (CLOCK_slo__sro_n50227));
AOI21_X2 CLOCK_slo__sro_c54928 (.ZN (CLOCK_slo__sro_n50224), .A (CLOCK_slo__sro_n50225)
    , .B1 (n_6_1520), .B2 (slo___n23247));
NAND2_X2 CLOCK_slo__sro_c55008 (.ZN (CLOCK_slo__sro_n50302), .A1 (n_6_859), .A2 (slo___n23463));
NAND2_X2 CLOCK_slo__sro_c55009 (.ZN (CLOCK_slo__sro_n50301), .A1 (CLOCK_slo__sro_n50302), .A2 (CLOCK_slo__sro_n50303));
AOI21_X2 CLOCK_slo__sro_c55010 (.ZN (CLOCK_slo__sro_n50300), .A (CLOCK_slo__sro_n50301)
    , .B1 (n_6_891), .B2 (slo___n23451));
INV_X2 CLOCK_slo__sro_c55026 (.ZN (CLOCK_slo__sro_n50320), .A (n_6_409));
BUF_X2 CLOCK_opt_ipo_c50602 (.Z (CLOCK_opt_ipo_n46265), .A (opt_ipo_n26244));
INV_X1 CLOCK_slo__sro_c55027 (.ZN (CLOCK_slo__sro_n50319), .A (n_6_1_904));
OAI21_X2 CLOCK_slo__sro_c55028 (.ZN (CLOCK_slo__sro_n50318), .A (CLOCK_slo__sro_n50321)
    , .B1 (CLOCK_slo__sro_n50320), .B2 (CLOCK_slo__sro_n50319));
AOI21_X4 CLOCK_slo__sro_c55029 (.ZN (slo__sro_n8965), .A (CLOCK_slo__sro_n50318), .B1 (n_6_441), .B2 (n_6_1_905));
NAND2_X1 CLOCK_slo__sro_c55042 (.ZN (CLOCK_slo__sro_n50331), .A1 (n_6_1_660), .A2 (n_6_866));
NAND2_X1 CLOCK_slo__sro_c55043 (.ZN (CLOCK_slo__sro_n50330), .A1 (CLOCK_slo__sro_n50331), .A2 (CLOCK_slo__sro_n50332));
AOI21_X4 CLOCK_slo__sro_c55044 (.ZN (slo__sro_n21560), .A (CLOCK_slo__sro_n50330)
    , .B1 (n_6_834), .B2 (slo___n23463));
NAND2_X1 CLOCK_slo__sro_c55078 (.ZN (CLOCK_slo__sro_n50363), .A1 (n_6_1_694), .A2 (n_6_782));
NAND2_X1 CLOCK_slo__sro_c55079 (.ZN (CLOCK_slo__sro_n50362), .A1 (CLOCK_slo__sro_n50363), .A2 (CLOCK_slo__sro_n50364));
AOI21_X1 CLOCK_slo__sro_c55080 (.ZN (n_6_1_675), .A (CLOCK_slo__sro_n50362), .B1 (n_6_814), .B2 (n_6_1_695));
NAND2_X1 CLOCK_slo__sro_c55122 (.ZN (CLOCK_slo__sro_n50402), .A1 (n_6_460), .A2 (n_6_1_869));
NAND2_X1 CLOCK_slo__sro_c55123 (.ZN (CLOCK_slo__sro_n50401), .A1 (CLOCK_slo__sro_n50402), .A2 (CLOCK_slo__sro_n50403));
AOI21_X2 CLOCK_slo__sro_c55124 (.ZN (CLOCK_slo__sro_n50400), .A (CLOCK_slo__sro_n50401)
    , .B1 (n_6_492), .B2 (n_6_1_870));
NAND2_X1 CLOCK_slo__sro_c55157 (.ZN (CLOCK_slo__sro_n50433), .A1 (n_6_967), .A2 (slo___n23232));
NAND2_X1 CLOCK_sgo__sro_c51309 (.ZN (CLOCK_sgo__sro_n47111), .A1 (n_6_2101), .A2 (n_6_1_168));
INV_X32 CLOCK_slo__c55145 (.ZN (n_6_1_274), .A (CLOCK_slo__n50421));
NAND2_X1 CLOCK_slo__sro_c55158 (.ZN (CLOCK_slo__sro_n50432), .A1 (CLOCK_slo__sro_n50433), .A2 (slo__sro_n40371));
INV_X2 CLOCK_slo__c59551 (.ZN (CLOCK_slo__n54206), .A (n_6_1_433));
NOR2_X2 CLOCK_slo__sro_c55216 (.ZN (slo__sro_n14081), .A1 (CLOCK_slo__sro_n50484), .A2 (slo__sro_n14082));
NAND2_X1 CLOCK_slo__sro_c55258 (.ZN (CLOCK_slo__sro_n50524), .A1 (slo___n23364), .A2 (n_6_1162));
NAND2_X1 CLOCK_slo__sro_c55259 (.ZN (CLOCK_slo__sro_n50523), .A1 (CLOCK_slo__sro_n50524), .A2 (CLOCK_slo__sro_n50525));
AOI21_X1 CLOCK_slo__sro_c55260 (.ZN (CLOCK_slo__sro_n50522), .A (CLOCK_slo__sro_n50523)
    , .B1 (n_6_1194), .B2 (slo___n23466));
AOI21_X2 CLOCK_slo__sro_c55353 (.ZN (CLOCK_slo__sro_n50608), .A (CLOCK_slo__sro_n50609)
    , .B1 (n_6_904), .B2 (slo___n23367));
AOI21_X2 CLOCK_slo__sro_c58617 (.ZN (n_6_1_444), .A (CLOCK_slo__sro_n53419), .B1 (n_6_1276), .B2 (slo___n23274));
NAND2_X1 CLOCK_slo__sro_c55350 (.ZN (CLOCK_slo__sro_n50611), .A1 (n_6_2488), .A2 (n_6_1_623));
NAND2_X2 CLOCK_slo__sro_c55351 (.ZN (CLOCK_slo__sro_n50610), .A1 (n_6_936), .A2 (n_6_1_625));
NAND2_X2 CLOCK_slo__sro_c55352 (.ZN (CLOCK_slo__sro_n50609), .A1 (CLOCK_slo__sro_n50610), .A2 (CLOCK_slo__sro_n50611));
NAND2_X1 CLOCK_slo__sro_c55402 (.ZN (CLOCK_slo__sro_n50658), .A1 (CLOCK_slo__sro_n50659), .A2 (CLOCK_slo__sro_n50660));
AOI21_X2 CLOCK_slo__sro_c55403 (.ZN (CLOCK_slo__sro_n50657), .A (CLOCK_slo__sro_n50658)
    , .B1 (n_6_1038), .B2 (n_6_1_554));
AOI222_X2 CLOCK_slo__sro_c72904 (.ZN (CLOCK_slo__n49050), .A1 (n_6_643), .A2 (n_6_1_764)
    , .B1 (n_6_675), .B2 (n_6_1_765), .C1 (n_6_2607), .C2 (n_6_1_763));
AND2_X1 CLOCK_slo__sro_c65721 (.ZN (CLOCK_slo__sro_n59232), .A1 (slo__sro_n7405), .A2 (n_6_1_518));
NOR2_X2 CLOCK_slo__sro_c55481 (.ZN (CLOCK_slo__sro_n50730), .A1 (CLOCK_slo__sro_n50731), .A2 (slo__sro_n15183));
NAND2_X1 CLOCK_slo__sro_c55543 (.ZN (CLOCK_slo__sro_n50793), .A1 (n_6_213), .A2 (n_6_1_1009));
NAND2_X1 CLOCK_slo__sro_c55544 (.ZN (CLOCK_slo__sro_n50792), .A1 (CLOCK_slo__sro_n50793), .A2 (CLOCK_slo__sro_n50794));
AOI21_X1 CLOCK_slo__sro_c55545 (.ZN (slo__sro_n13965), .A (CLOCK_slo__sro_n50792)
    , .B1 (n_6_245), .B2 (n_6_1_1010));
NAND2_X1 CLOCK_slo__sro_c55588 (.ZN (CLOCK_slo__sro_n50831), .A1 (n_6_141), .A2 (n_6_1_1044));
NAND2_X1 CLOCK_slo__sro_c55589 (.ZN (CLOCK_slo__sro_n50830), .A1 (CLOCK_slo__sro_n50831), .A2 (slo__sro_n20974));
AOI21_X1 CLOCK_slo__sro_c55590 (.ZN (n_6_1_1024), .A (CLOCK_slo__sro_n50830), .B1 (n_6_173), .B2 (n_6_1_1045));
INV_X1 CLOCK_slo__sro_c55602 (.ZN (CLOCK_slo__sro_n50840), .A (CLOCK_slo__sro_n50841));
NOR2_X1 CLOCK_slo__sro_c55603 (.ZN (slo__sro_n29674), .A1 (slo__sro_n29675), .A2 (CLOCK_slo__sro_n50840));
NOR2_X2 CLOCK_slo__sro_c55616 (.ZN (slo__sro_n32470), .A1 (CLOCK_slo__sro_n50850), .A2 (slo__sro_n32471));
NAND2_X1 CLOCK_slo__sro_c55632 (.ZN (CLOCK_slo__sro_n50863), .A1 (n_6_267), .A2 (n_6_1_974));
NAND2_X1 CLOCK_slo__sro_c55633 (.ZN (CLOCK_slo__sro_n50862), .A1 (CLOCK_slo__sro_n50863), .A2 (CLOCK_slo__sro_n50864));
AOI21_X1 CLOCK_slo__sro_c55634 (.ZN (slo__sro_n10838), .A (CLOCK_slo__sro_n50862)
    , .B1 (n_6_299), .B2 (n_6_1_975));
AOI21_X1 CLOCK_slo__sro_c55689 (.ZN (CLOCK_slo__sro_n50912), .A (slo__sro_n19998)
    , .B1 (n_6_1226), .B2 (slo___n23359));
AND2_X1 CLOCK_slo__sro_c55690 (.ZN (slo__sro_n19997), .A1 (CLOCK_slo__sro_n50913), .A2 (CLOCK_slo__sro_n50912));
NAND2_X1 CLOCK_slo__sro_c55755 (.ZN (CLOCK_slo__sro_n50975), .A1 (n_6_686), .A2 (n_6_1_765));
NAND2_X1 CLOCK_slo__sro_c55756 (.ZN (CLOCK_slo__sro_n50974), .A1 (CLOCK_slo__sro_n50975), .A2 (CLOCK_slo__sro_n50976));
AOI21_X1 CLOCK_slo__sro_c55757 (.ZN (n_6_1_745), .A (CLOCK_slo__sro_n50974), .B1 (n_6_654), .B2 (n_6_1_764));
AOI21_X1 CLOCK_slo__sro_c55774 (.ZN (CLOCK_slo__sro_n50986), .A (slo__sro_n7038), .B1 (n_6_1500), .B2 (n_6_1_309));
AND2_X1 CLOCK_slo__sro_c55775 (.ZN (slo__sro_n7037), .A1 (CLOCK_slo__sro_n50987), .A2 (CLOCK_slo__sro_n50986));
AOI21_X2 CLOCK_slo__sro_c55857 (.ZN (CLOCK_slo__sro_n51061), .A (slo__sro_n7098), .B1 (n_6_1492), .B2 (n_6_1_309));
AND2_X1 CLOCK_slo__sro_c55858 (.ZN (CLOCK_slo__sro_n51060), .A1 (CLOCK_slo__sro_n51061), .A2 (CLOCK_slo__sro_n51062));
NAND2_X1 CLOCK_slo__sro_c55892 (.ZN (CLOCK_slo__sro_n51094), .A1 (n_6_1_764), .A2 (n_6_656));
NAND2_X1 CLOCK_slo__sro_c55893 (.ZN (CLOCK_slo__sro_n51093), .A1 (CLOCK_slo__sro_n51094), .A2 (CLOCK_slo__sro_n51095));
AOI21_X2 CLOCK_slo__sro_c55894 (.ZN (CLOCK_slo__sro_n51092), .A (CLOCK_slo__sro_n51093)
    , .B1 (n_6_688), .B2 (n_6_1_765));
AOI221_X2 CLOCK_slo__sro_c55933 (.ZN (CLOCK_slo__sro_n51132), .A (CLOCK_slo__sro_n51133)
    , .B1 (n_6_997), .B2 (slo___n23218), .C1 (n_6_965), .C2 (slo___n23232));
INV_X2 CLOCK_slo__c55997 (.ZN (slo__sro_n30921), .A (CLOCK_slo__sro_n53156));
NAND2_X1 CLOCK_slo__sro_c56072 (.ZN (CLOCK_slo__sro_n51260), .A1 (CLOCK_slo__sro_n51261), .A2 (CLOCK_slo__sro_n51262));
AOI21_X2 CLOCK_slo__sro_c56073 (.ZN (n_6_1_793), .A (CLOCK_slo__sro_n51260), .B1 (n_6_635), .B2 (n_6_1_800));
INV_X2 opt_ipo_c48942 (.ZN (opt_ipo_n44599), .A (slo__sro_n35249));
NAND2_X1 CLOCK_slo__sro_c56122 (.ZN (CLOCK_slo__sro_n51307), .A1 (CLOCK_slo__sro_n51309), .A2 (CLOCK_slo__sro_n51308));
AOI21_X1 CLOCK_slo__sro_c56123 (.ZN (CLOCK_slo__sro_n51306), .A (CLOCK_slo__sro_n51307)
    , .B1 (n_6_174), .B2 (n_6_1_1045));
NAND2_X2 CLOCK_slo__mro_c56197 (.ZN (CLOCK_slo__mro_n51373), .A1 (n_6_1436), .A2 (slo___n23229));
NAND2_X2 CLOCK_slo__mro_c56198 (.ZN (CLOCK_slo__mro_n51372), .A1 (CLOCK_slo__mro_n51373), .A2 (slo__sro_n9794));
NOR2_X4 CLOCK_slo__mro_c56199 (.ZN (CLOCK_slo__mro_n51371), .A1 (CLOCK_slo__mro_n51372), .A2 (slo__sro_n39872));
AOI21_X2 CLOCK_slo__sro_c56311 (.ZN (n_6_1_201), .A (CLOCK_slo__sro_n51473), .B1 (n_6_1726), .B2 (slo___n23407));
NAND2_X1 CLOCK_slo__sro_c56274 (.ZN (CLOCK_slo__sro_n51442), .A1 (n_6_1_623), .A2 (n_6_2499));
NAND2_X1 CLOCK_slo__sro_c56275 (.ZN (CLOCK_slo__sro_n51441), .A1 (n_6_915), .A2 (slo___n23367));
NAND2_X1 CLOCK_slo__sro_c56276 (.ZN (CLOCK_slo__sro_n51440), .A1 (CLOCK_slo__sro_n51441), .A2 (CLOCK_slo__sro_n51442));
AOI21_X1 CLOCK_slo__sro_c56277 (.ZN (CLOCK_slo__sro_n51439), .A (CLOCK_slo__sro_n51440)
    , .B1 (n_6_947), .B2 (n_6_1_625));
NAND2_X1 CLOCK_slo__mro_c56342 (.ZN (CLOCK_slo__mro_n51497), .A1 (n_6_998), .A2 (slo___n23218));
NAND2_X1 CLOCK_slo__mro_c56343 (.ZN (slo__sro_n17951), .A1 (CLOCK_slo__mro_n51497), .A2 (slo__sro_n17953));
INV_X1 CLOCK_slo__mro_c56381 (.ZN (CLOCK_slo__mro_n51529), .A (slo___n23274));
INV_X1 CLOCK_slo__mro_c56382 (.ZN (slo__sro_n19545), .A (n_6_1254));
OAI21_X1 CLOCK_slo__mro_c56383 (.ZN (slo__sro_n19544), .A (slo__sro_n19546), .B1 (slo__sro_n19545), .B2 (CLOCK_slo__mro_n51529));
AOI221_X2 CLOCK_slo__sro_c56462 (.ZN (slo__sro_n15534), .A (CLOCK_slo__sro_n51595)
    , .B1 (n_6_1771), .B2 (CLOCK_sgo__n48020), .C1 (n_6_1739), .C2 (n_6_1_169));
NAND2_X1 CLOCK_slo__sro_c56472 (.ZN (CLOCK_slo__sro_n51603), .A1 (n_6_1605), .A2 (slo___n23215));
NAND2_X1 CLOCK_slo__sro_c56473 (.ZN (CLOCK_slo__sro_n51602), .A1 (CLOCK_slo__sro_n51603), .A2 (CLOCK_slo__sro_n51604));
AOI21_X2 CLOCK_slo__sro_c56474 (.ZN (CLOCK_slo__sro_n51601), .A (CLOCK_slo__sro_n51602)
    , .B1 (n_6_1637), .B2 (drc_ipo_n26601));
NAND2_X1 CLOCK_slo__sro_c56490 (.ZN (CLOCK_slo__sro_n51620), .A1 (n_6_1_869), .A2 (n_6_461));
NAND2_X1 CLOCK_slo__sro_c56491 (.ZN (CLOCK_slo__sro_n51619), .A1 (CLOCK_slo__sro_n51620), .A2 (CLOCK_slo__sro_n51621));
NAND2_X1 CLOCK_slo__sro_c71928 (.ZN (CLOCK_slo__sro_n64637), .A1 (CLOCK_slo__sro_n64639), .A2 (CLOCK_slo__sro_n64638));
NAND2_X1 CLOCK_slo__sro_c56518 (.ZN (CLOCK_slo__sro_n51645), .A1 (n_6_1_835), .A2 (n_6_559));
NAND2_X1 CLOCK_slo__sro_c56519 (.ZN (CLOCK_slo__sro_n51644), .A1 (CLOCK_slo__sro_n51645), .A2 (slo__sro_n5270));
AOI21_X1 CLOCK_slo__sro_c56520 (.ZN (CLOCK_slo__sro_n51643), .A (CLOCK_slo__sro_n51644)
    , .B1 (n_6_527), .B2 (n_6_1_834));
AOI21_X1 CLOCK_slo__sro_c56613 (.ZN (CLOCK_slo__sro_n51724), .A (slo__sro_n15199)
    , .B1 (n_6_623), .B2 (n_6_1_800));
NAND2_X1 CLOCK_sgo__sro_c51478 (.ZN (CLOCK_sgo__sro_n47244), .A1 (CLOCK_sgo__sro_n47245), .A2 (CLOCK_sgo__sro_n47246));
AND2_X2 CLOCK_slo__sro_c56614 (.ZN (CLOCK_slo__sro_n51723), .A1 (CLOCK_slo__sro_n51724), .A2 (CLOCK_slo__sro_n51725));
AOI21_X1 CLOCK_slo__sro_c56662 (.ZN (CLOCK_slo__sro_n51765), .A (n_6_1_692), .B1 (n_6_797), .B2 (n_6_1_694));
AND2_X1 CLOCK_slo__sro_c56663 (.ZN (n_6_1_690), .A1 (CLOCK_slo__sro_n51765), .A2 (CLOCK_slo__sro_n51766));
NAND2_X1 CLOCK_slo__sro_c56675 (.ZN (CLOCK_slo__sro_n51774), .A1 (CLOCK_slo__sro_n51775), .A2 (CLOCK_slo__sro_n51776));
AOI21_X1 CLOCK_slo__sro_c56676 (.ZN (CLOCK_slo__sro_n51773), .A (CLOCK_slo__sro_n51774)
    , .B1 (n_6_1870), .B2 (CLOCK_sgo__n48011));
INV_X1 CLOCK_slo__sro_c56763 (.ZN (CLOCK_slo__sro_n51852), .A (CLOCK_slo__sro_n51853));
NAND2_X1 CLOCK_slo__sro_c59645 (.ZN (CLOCK_slo__sro_n54282), .A1 (CLOCK_sgo__n48020), .A2 (n_6_1780));
NOR2_X2 CLOCK_slo__sro_c56764 (.ZN (n_6_1_245), .A1 (slo__sro_n18154), .A2 (CLOCK_slo__sro_n51852));
INV_X1 CLOCK_slo__sro_c56800 (.ZN (CLOCK_slo__sro_n51886), .A (CLOCK_slo__sro_n51887));
NOR2_X4 CLOCK_slo__sro_c56801 (.ZN (CLOCK_slo__sro_n51885), .A1 (CLOCK_slo__sro_n51886), .A2 (slo__sro_n34756));
INV_X1 CLOCK_slo__sro_c56740 (.ZN (CLOCK_slo__sro_n51836), .A (n_6_1_587));
NAND2_X1 CLOCK_slo__sro_c56741 (.ZN (CLOCK_slo__sro_n51835), .A1 (n_6_1021), .A2 (slo___n23218));
NAND2_X1 CLOCK_slo__sro_c56742 (.ZN (CLOCK_slo__sro_n51834), .A1 (n_6_989), .A2 (slo___n23232));
AND3_X1 CLOCK_slo__sro_c56743 (.ZN (n_6_1_585), .A1 (CLOCK_slo__sro_n51835), .A2 (CLOCK_slo__sro_n51834), .A3 (CLOCK_slo__sro_n51836));
AND2_X1 CLOCK_slo__sro_c56907 (.ZN (CLOCK_slo__sro_n51957), .A1 (CLOCK_slo__sro_n51959), .A2 (CLOCK_slo__sro_n51958));
NAND2_X1 CLOCK_slo__sro_c56939 (.ZN (CLOCK_slo__sro_n51981), .A1 (n_6_1104), .A2 (slo___n23277));
NAND2_X2 CLOCK_slo__mro_c56918 (.ZN (slo__sro_n20323), .A1 (n_6_1100), .A2 (slo___n23277));
NAND2_X2 CLOCK_slo__mro_c56919 (.ZN (slo__sro_n20322), .A1 (slo__sro_n20323), .A2 (slo__sro_n20324));
NOR2_X1 CLOCK_slo__sro_c56968 (.ZN (slo__n39180), .A1 (slo__sro_n29489), .A2 (CLOCK_slo__sro_n52005));
INV_X1 CLOCK_slo__sro_c57130 (.ZN (CLOCK_slo__sro_n52125), .A (CLOCK_slo__sro_n52126));
NAND2_X1 CLOCK_slo__sro_c57681 (.ZN (CLOCK_slo__sro_n52595), .A1 (n_6_1_238), .A2 (n_6_2152));
INV_X1 CLOCK_slo__sro_c57142 (.ZN (CLOCK_slo__sro_n52137), .A (CLOCK_slo__sro_n52138));
NAND2_X1 CLOCK_slo__sro_c57024 (.ZN (CLOCK_slo__sro_n52056), .A1 (CLOCK_sgo__n46950), .A2 (n_6_2830));
NAND2_X1 CLOCK_slo__sro_c57025 (.ZN (CLOCK_slo__sro_n52055), .A1 (n_6_233), .A2 (n_6_1_1010));
NAND2_X1 CLOCK_slo__sro_c57026 (.ZN (CLOCK_slo__sro_n52054), .A1 (CLOCK_slo__sro_n52055), .A2 (CLOCK_slo__sro_n52056));
AOI21_X1 CLOCK_slo__sro_c57027 (.ZN (n_6_1_985), .A (CLOCK_slo__sro_n52054), .B1 (n_6_201), .B2 (n_6_1_1009));
AOI222_X2 CLOCK_slo__sro_c57231 (.ZN (slo__sro_n18343), .A1 (n_6_1281), .A2 (n_6_1_414)
    , .B1 (n_6_1313), .B2 (slo___n43257), .C1 (n_6_2295), .C2 (n_6_1_413));
INV_X2 CLOCK_slo__mro_c57175 (.ZN (CLOCK_slo__mro_n52164), .A (n_6_1559));
INV_X1 CLOCK_slo__mro_c57176 (.ZN (slo__sro_n15686), .A (CLOCK_sgo__n48008));
OAI21_X2 CLOCK_slo__mro_c57177 (.ZN (slo__sro_n15685), .A (slo__sro_n15687), .B1 (CLOCK_slo__mro_n52164), .B2 (slo__sro_n15686));
OAI21_X2 CLOCK_slo__mro_c57200 (.ZN (CLOCK_slo__mro_n52173), .A (slo__sro_n20568)
    , .B1 (CLOCK_slo__mro_n52174), .B2 (slo__sro_n42343));
NAND2_X1 CLOCK_slo__sro_c57682 (.ZN (CLOCK_slo__sro_n52594), .A1 (drc_ipo_n26601), .A2 (n_6_1645));
NAND2_X1 CLOCK_slo__sro_c57657 (.ZN (CLOCK_slo__sro_n52571), .A1 (n_6_2893), .A2 (slo__n13799));
NAND2_X1 CLOCK_slo__sro_c57658 (.ZN (CLOCK_slo__sro_n52570), .A1 (n_6_106), .A2 (n_6_1_1080));
AOI222_X2 CLOCK_slo__sro_c57272 (.ZN (n_6_1_630), .A1 (n_6_868), .A2 (n_6_1_660), .B1 (n_6_836)
    , .B2 (slo___n23463), .C1 (slo___n16283), .C2 (n_6_1_658));
AOI21_X1 CLOCK_slo__sro_c57660 (.ZN (CLOCK_slo__sro_n52568), .A (CLOCK_slo__sro_n52569)
    , .B1 (n_6_74), .B2 (n_6_1_1079));
NAND2_X1 CLOCK_slo__sro_c57625 (.ZN (CLOCK_slo__sro_n52542), .A1 (n_6_2266), .A2 (n_6_1_378));
NAND2_X1 CLOCK_slo__sro_c57626 (.ZN (CLOCK_slo__sro_n52541), .A1 (n_6_1347), .A2 (n_6_1_379));
NAND2_X1 CLOCK_slo__sro_c57627 (.ZN (CLOCK_slo__sro_n52540), .A1 (CLOCK_slo__sro_n52541), .A2 (CLOCK_slo__sro_n52542));
AOI21_X2 CLOCK_slo__sro_c57628 (.ZN (n_6_1_349), .A (CLOCK_slo__sro_n52540), .B1 (n_6_1379), .B2 (n_6_1_380));
NAND2_X1 CLOCK_slo__sro_c57760 (.ZN (CLOCK_slo__sro_n52669), .A1 (CLOCK_slo__sro_n52670), .A2 (CLOCK_slo__sro_n52671));
AOI21_X2 CLOCK_slo__sro_c57761 (.ZN (slo__sro_n33384), .A (CLOCK_slo__sro_n52669)
    , .B1 (n_6_1014), .B2 (slo___n23218));
INV_X1 CLOCK_slo__sro_c57721 (.ZN (CLOCK_slo__sro_n52635), .A (slo__sro_n9916));
NAND2_X1 CLOCK_slo__sro_c57722 (.ZN (CLOCK_slo__sro_n52634), .A1 (n_6_1372), .A2 (n_6_1_379));
NAND2_X1 CLOCK_slo__sro_c57723 (.ZN (CLOCK_slo__sro_n52633), .A1 (CLOCK_slo__sro_n52634), .A2 (CLOCK_slo__sro_n52635));
AOI21_X2 CLOCK_slo__sro_c58033 (.ZN (n_6_1_166), .A (CLOCK_slo__sro_n52915), .B1 (n_6_1790), .B2 (n_6_1_170));
NAND2_X1 CLOCK_slo__sro_c58102 (.ZN (CLOCK_slo__sro_n52972), .A1 (n_6_217), .A2 (n_6_1_1009));
AOI21_X2 CLOCK_slo__sro_c57724 (.ZN (CLOCK_slo__sro_n52632), .A (CLOCK_slo__sro_n52633)
    , .B1 (n_6_1404), .B2 (n_6_1_380));
AOI222_X2 CLOCK_slo__sro_c57539 (.ZN (CLOCK_slo__sro_n52466), .A1 (n_6_1235), .A2 (slo___n23359)
    , .B1 (n_6_1267), .B2 (slo___n23274), .C1 (n_6_2344), .C2 (n_6_1_448));
AOI21_X1 CLOCK_slo__sro_c58103 (.ZN (CLOCK_slo__sro_n52971), .A (slo__sro_n22623)
    , .B1 (n_6_249), .B2 (n_6_1_1010));
AND2_X1 CLOCK_slo__sro_c58104 (.ZN (n_6_1_1001), .A1 (CLOCK_slo__sro_n52972), .A2 (CLOCK_slo__sro_n52971));
NAND2_X1 CLOCK_slo__sro_c58225 (.ZN (CLOCK_slo__sro_n53079), .A1 (n_6_105), .A2 (n_6_1_1080));
NAND2_X1 CLOCK_slo__sro_c58226 (.ZN (CLOCK_slo__sro_n53078), .A1 (CLOCK_slo__sro_n53080), .A2 (CLOCK_slo__sro_n53079));
AOI222_X2 CLOCK_slo__sro_c58153 (.ZN (CLOCK_slo__sro_n53015), .A1 (n_6_555), .A2 (n_6_1_835)
    , .B1 (n_6_523), .B2 (n_6_1_834), .C1 (CLOCK_slo__n58182), .C2 (CLOCK_sgo__n46922));
NAND2_X1 CLOCK_slo__sro_c57897 (.ZN (CLOCK_slo__sro_n52795), .A1 (n_6_1_274), .A2 (n_6_1548));
NAND2_X1 CLOCK_slo__sro_c57898 (.ZN (CLOCK_slo__sro_n52794), .A1 (CLOCK_slo__sro_n52795), .A2 (slo__sro_n38324));
AOI21_X2 CLOCK_slo__sro_c57899 (.ZN (slo__n28105), .A (CLOCK_slo__sro_n52794), .B1 (n_6_1580), .B2 (slo___n23244));
AOI222_X2 CLOCK_slo__sro_c58288 (.ZN (n_6_1_252), .A1 (n_6_1579), .A2 (slo___n23244)
    , .B1 (n_6_1547), .B2 (n_6_1_274), .C1 (n_6_2181), .C2 (n_6_1_273));
NAND2_X1 CLOCK_slo__sro_c58455 (.ZN (CLOCK_slo__sro_n53278), .A1 (n_6_1_274), .A2 (n_6_1564));
AND2_X1 CLOCK_slo__sro_c58206 (.ZN (CLOCK_slo__sro_n53064), .A1 (n_6_2659), .A2 (n_6_1_798));
AOI221_X2 CLOCK_slo__sro_c58207 (.ZN (n_6_1_790), .A (CLOCK_slo__sro_n53064), .B1 (n_6_600)
    , .B2 (n_6_1_799), .C1 (n_6_632), .C2 (n_6_1_800));
NAND2_X1 CLOCK_slo__sro_c58325 (.ZN (CLOCK_slo__sro_n53158), .A1 (slo___n23239), .A2 (n_6_1672));
NAND2_X1 CLOCK_slo__sro_c58326 (.ZN (CLOCK_slo__sro_n53157), .A1 (CLOCK_slo__sro_n53158), .A2 (CLOCK_slo__sro_n53159));
AOI21_X1 CLOCK_slo__sro_c58327 (.ZN (CLOCK_slo__sro_n53156), .A (CLOCK_slo__sro_n53157)
    , .B1 (n_6_1704), .B2 (slo___n23407));
INV_X2 CLOCK_slo__c58684 (.ZN (CLOCK_slo__n53479), .A (n_6_1_329));
NAND2_X1 CLOCK_slo__sro_c58364 (.ZN (CLOCK_slo__sro_n53198), .A1 (n_6_2283), .A2 (n_6_1_378));
INV_X1 CLOCK_slo__sro_c58365 (.ZN (CLOCK_slo__sro_n53197), .A (CLOCK_slo__sro_n53198));
AOI221_X2 CLOCK_slo__sro_c58366 (.ZN (CLOCK_slo__sro_n53196), .A (CLOCK_slo__sro_n53197)
    , .B1 (n_6_1364), .B2 (n_6_1_379), .C1 (n_6_1396), .C2 (n_6_1_380));
NAND2_X1 CLOCK_slo__sro_c58597 (.ZN (CLOCK_slo__sro_n53406), .A1 (n_6_1039), .A2 (n_6_1_554));
NAND2_X1 CLOCK_slo__sro_c58598 (.ZN (CLOCK_slo__sro_n53405), .A1 (CLOCK_slo__sro_n53406), .A2 (CLOCK_slo__sro_n50547));
AOI21_X1 CLOCK_slo__sro_c58599 (.ZN (n_6_1_536), .A (CLOCK_slo__sro_n53405), .B1 (n_6_1071), .B2 (slo___n23457));
INV_X1 CLOCK_slo__sro_c58792 (.ZN (CLOCK_slo__sro_n53571), .A (CLOCK_slo__sro_n53572));
INV_X1 CLOCK_slo__sro_c58431 (.ZN (CLOCK_slo__sro_n53260), .A (slo__sro_n23125));
NAND2_X1 CLOCK_slo__sro_c58432 (.ZN (CLOCK_slo__sro_n53259), .A1 (n_6_1416), .A2 (slo___n23229));
NAND2_X2 CLOCK_slo__sro_c58433 (.ZN (CLOCK_slo__sro_n53258), .A1 (CLOCK_slo__sro_n53259), .A2 (CLOCK_slo__sro_n53260));
AOI21_X4 CLOCK_slo__sro_c58434 (.ZN (CLOCK_slo__sro_n53257), .A (CLOCK_slo__sro_n53258)
    , .B1 (n_6_1448), .B2 (n_6_1_345));
AOI221_X2 CLOCK_slo__sro_c58793 (.ZN (n_6_1_217), .A (CLOCK_slo__sro_n53571), .B1 (n_6_1643)
    , .B2 (drc_ipo_n26601), .C1 (n_6_1611), .C2 (slo___n23215));
AOI222_X2 CLOCK_slo__sro_c71299 (.ZN (n_6_1_572), .A1 (n_6_976), .A2 (slo___n23232)
    , .B1 (n_6_1008), .B2 (slo___n23218), .C1 (n_6_2465), .C2 (n_6_1_588));
NAND2_X1 CLOCK_slo__sro_c59682 (.ZN (CLOCK_slo__sro_n54315), .A1 (n_6_2053), .A2 (n_6_1_133));
INV_X1 CLOCK_slo__c58960 (.ZN (CLOCK_slo__n53697), .A (slo__sro_n7557));
NAND2_X1 CLOCK_slo__sro_c59416 (.ZN (CLOCK_slo__sro_n54101), .A1 (drc_ipo_n26601), .A2 (n_6_1656));
INV_X1 CLOCK_slo__sro_c59370 (.ZN (CLOCK_slo__sro_n54056), .A (slo__sro_n5711));
NAND2_X1 CLOCK_slo__sro_c59371 (.ZN (CLOCK_slo__sro_n54055), .A1 (n_6_1072), .A2 (slo___n23457));
NAND2_X1 CLOCK_slo__sro_c59102 (.ZN (CLOCK_slo__sro_n53825), .A1 (n_6_2205), .A2 (n_6_1_308));
NAND2_X1 CLOCK_slo__sro_c59103 (.ZN (CLOCK_slo__sro_n53824), .A1 (n_6_1_309), .A2 (n_6_1476));
NAND2_X1 CLOCK_slo__sro_c59104 (.ZN (CLOCK_slo__sro_n53823), .A1 (CLOCK_slo__sro_n53824), .A2 (CLOCK_slo__sro_n53825));
AOI21_X2 CLOCK_slo__sro_c59105 (.ZN (n_6_1_280), .A (CLOCK_slo__sro_n53823), .B1 (n_6_1508), .B2 (slo___n23247));
AND3_X1 CLOCK_slo__sro_c59373 (.ZN (CLOCK_slo__sro_n54053), .A1 (CLOCK_slo__sro_n54054)
    , .A2 (CLOCK_slo__sro_n54056), .A3 (CLOCK_slo__sro_n54055));
NAND2_X1 CLOCK_slo__sro_c59220 (.ZN (CLOCK_slo__sro_n53932), .A1 (n_6_999), .A2 (slo___n23218));
NAND2_X1 CLOCK_slo__sro_c59175 (.ZN (CLOCK_slo__sro_n53894), .A1 (n_6_1341), .A2 (slo___n43257));
AOI21_X1 CLOCK_slo__sro_c59176 (.ZN (CLOCK_slo__sro_n53893), .A (n_6_1_412), .B1 (n_6_1309), .B2 (n_6_1_414));
AND2_X1 CLOCK_slo__sro_c59177 (.ZN (CLOCK_slo__sro_n53892), .A1 (CLOCK_slo__sro_n53894), .A2 (CLOCK_slo__sro_n53893));
NOR2_X2 CLOCK_slo__sro_c59222 (.ZN (n_6_1_563), .A1 (CLOCK_slo__sro_n50432), .A2 (CLOCK_slo__sro_n53931));
INV_X1 CLOCK_slo__c59529 (.ZN (CLOCK_slo__n54187), .A (CLOCK_slo__sro_n64180));
AOI222_X2 CLOCK_slo__sro_c59491 (.ZN (slo__sro_n14441), .A1 (n_6_1674), .A2 (slo___n23239)
    , .B1 (n_6_1706), .B2 (slo___n23407), .C1 (opt_ipo_n24541), .C2 (n_6_1_203));
AOI21_X1 CLOCK_slo__sro_c59685 (.ZN (CLOCK_slo__sro_n54312), .A (CLOCK_slo__sro_n54313)
    , .B1 (n_6_1799), .B2 (n_6_1_134));
NAND2_X2 CLOCK_slo__sro_c59646 (.ZN (CLOCK_slo__sro_n54281), .A1 (CLOCK_slo__sro_n54282), .A2 (slo__sro_n27140));
AOI21_X2 CLOCK_slo__sro_c59647 (.ZN (slo__sro_n27138), .A (CLOCK_slo__sro_n54281)
    , .B1 (n_6_1748), .B2 (n_6_1_169));
NAND2_X1 CLOCK_slo__sro_c59683 (.ZN (CLOCK_slo__sro_n54314), .A1 (n_6_1831), .A2 (n_6_1_135));
NAND2_X1 CLOCK_slo__sro_c59684 (.ZN (CLOCK_slo__sro_n54313), .A1 (CLOCK_slo__sro_n54314), .A2 (CLOCK_slo__sro_n54315));
INV_X1 CLOCK_slo__sro_c59890 (.ZN (CLOCK_slo__sro_n54488), .A (CLOCK_slo__sro_n54489));
NAND2_X1 CLOCK_slo__sro_c59873 (.ZN (CLOCK_slo__sro_n54474), .A1 (n_6_2114), .A2 (n_6_1_203));
NAND2_X1 CLOCK_slo__sro_c59874 (.ZN (CLOCK_slo__sro_n54473), .A1 (n_6_1670), .A2 (slo___n23239));
NAND2_X1 CLOCK_slo__sro_c59875 (.ZN (CLOCK_slo__sro_n54472), .A1 (CLOCK_slo__sro_n54474), .A2 (CLOCK_slo__sro_n54473));
AOI21_X1 CLOCK_slo__sro_c59876 (.ZN (CLOCK_slo__sro_n54471), .A (CLOCK_slo__sro_n54472)
    , .B1 (n_6_1702), .B2 (slo___n23407));
NAND2_X1 CLOCK_slo__sro_c59976 (.ZN (CLOCK_slo__sro_n54568), .A1 (n_6_1512), .A2 (slo___n23247));
NAND2_X1 CLOCK_slo__sro_c59977 (.ZN (CLOCK_slo__sro_n54567), .A1 (n_6_1480), .A2 (n_6_1_309));
AND3_X1 CLOCK_slo__sro_c59978 (.ZN (slo__sro_n29225), .A1 (CLOCK_slo__sro_n54568)
    , .A2 (CLOCK_slo__sro_n54569), .A3 (CLOCK_slo__sro_n54567));
AND2_X1 CLOCK_slo__sro_c60024 (.ZN (CLOCK_slo__sro_n54605), .A1 (n_6_1315), .A2 (slo___n43257));
NOR2_X2 CLOCK_slo__sro_c60025 (.ZN (n_6_1_384), .A1 (slo__sro_n6689), .A2 (CLOCK_slo__sro_n54605));
AOI222_X2 CLOCK_slo__sro_c60076 (.ZN (CLOCK_slo__sro_n54647), .A1 (n_6_745), .A2 (n_6_1_730)
    , .B1 (n_6_713), .B2 (n_6_1_729), .C1 (n_6_2582), .C2 (n_6_1_728));
NOR2_X4 CLOCK_slo__sro_c60134 (.ZN (n_6_1_969), .A1 (CLOCK_slo__sro_n54698), .A2 (slo__sro_n31670));
INV_X1 CLOCK_slo__sro_c59959 (.ZN (CLOCK_slo__sro_n54554), .A (n_6_2561));
INV_X1 CLOCK_slo__sro_c59960 (.ZN (CLOCK_slo__sro_n54553), .A (n_6_1_693));
NOR2_X1 CLOCK_slo__sro_c59961 (.ZN (CLOCK_slo__sro_n54552), .A1 (CLOCK_slo__sro_n54554), .A2 (CLOCK_slo__sro_n54553));
AOI221_X2 CLOCK_slo__sro_c59962 (.ZN (CLOCK_slo__sro_n54551), .A (CLOCK_slo__sro_n54552)
    , .B1 (n_6_787), .B2 (n_6_1_694), .C1 (n_6_819), .C2 (n_6_1_695));
AOI221_X2 CLOCK_slo__sro_c60147 (.ZN (n_6_1_103), .A (CLOCK_slo__sro_n54706), .B1 (n_6_1794)
    , .B2 (n_6_1_134), .C1 (n_6_1826), .C2 (slo___n23404));
AOI21_X1 CLOCK_slo__sro_c69833 (.ZN (slo__sro_n40769), .A (CLOCK_slo__sro_n62893)
    , .B1 (n_6_188), .B2 (n_6_1_1045));
NAND2_X1 CLOCK_slo__sro_c60343 (.ZN (CLOCK_slo__sro_n54886), .A1 (n_6_524), .A2 (n_6_1_834));
NAND2_X1 CLOCK_slo__sro_c60344 (.ZN (CLOCK_slo__sro_n54885), .A1 (n_6_556), .A2 (n_6_1_835));
NAND3_X1 CLOCK_slo__sro_c60345 (.ZN (CLOCK_slo__sro_n54884), .A1 (CLOCK_slo__sro_n54885)
    , .A2 (CLOCK_slo__sro_n54886), .A3 (slo__sro_n5285));
INV_X1 CLOCK_slo__sro_c60346 (.ZN (n_6_1_813), .A (CLOCK_slo__sro_n54884));
AOI222_X2 CLOCK_slo__sro_c60235 (.ZN (CLOCK_slo__sro_n54789), .A1 (n_6_1810), .A2 (n_6_1_134)
    , .B1 (n_6_1842), .B2 (n_6_1_135), .C1 (n_6_2064), .C2 (n_6_1_133));
INV_X2 CLOCK_slo__c60541 (.ZN (slo__sro_n7405), .A (CLOCK_slo__n55041));
NOR2_X1 CLOCK_slo__sro_c60560 (.ZN (CLOCK_slo__sro_n55059), .A1 (slo__sro_n40148), .A2 (CLOCK_slo__sro_n55060));
OAI21_X1 CLOCK_slo__sro_c60519 (.ZN (CLOCK_slo__sro_n55020), .A (CLOCK_slo__sro_n55023)
    , .B1 (CLOCK_slo__sro_n55022), .B2 (CLOCK_slo__sro_n55021));
AND2_X1 CLOCK_slo__sro_c60429 (.ZN (CLOCK_slo__sro_n54952), .A1 (n_6_88), .A2 (n_6_1_1079));
NOR2_X1 CLOCK_slo__sro_c60430 (.ZN (slo__sro_n7944), .A1 (slo__sro_n7945), .A2 (CLOCK_slo__sro_n54952));
AOI21_X2 CLOCK_slo__sro_c60520 (.ZN (CLOCK_slo__sro_n55019), .A (CLOCK_slo__sro_n55020)
    , .B1 (n_6_1269), .B2 (slo___n23274));
INV_X2 CLOCK_slo__c60579 (.ZN (CLOCK_slo__n55073), .A (slo__sro_n41478));
AOI222_X2 CLOCK_slo__sro_c60494 (.ZN (n_6_1_557), .A1 (n_6_993), .A2 (slo___n23218)
    , .B1 (n_6_961), .B2 (slo___n23232), .C1 (n_6_2450), .C2 (n_6_1_588));
NAND2_X1 CLOCK_slo__sro_c60595 (.ZN (CLOCK_slo__sro_n55085), .A1 (CLOCK_slo__sro_n55086), .A2 (CLOCK_slo__sro_n55087));
AOI21_X1 CLOCK_slo__sro_c60596 (.ZN (CLOCK_slo__sro_n55084), .A (CLOCK_slo__sro_n55085)
    , .B1 (n_6_1444), .B2 (n_6_1_345));
INV_X1 CLOCK_slo__sro_c60612 (.ZN (CLOCK_slo__sro_n55104), .A (n_6_1_693));
NOR2_X1 CLOCK_slo__sro_c60613 (.ZN (CLOCK_slo__sro_n55103), .A1 (CLOCK_slo__sro_n55105), .A2 (CLOCK_slo__sro_n55104));
AOI221_X2 CLOCK_slo__sro_c60614 (.ZN (CLOCK_slo__sro_n55102), .A (CLOCK_slo__sro_n55103)
    , .B1 (n_6_796), .B2 (n_6_1_694), .C1 (n_6_828), .C2 (n_6_1_695));
NAND2_X1 CLOCK_slo__sro_c60697 (.ZN (CLOCK_slo__sro_n55170), .A1 (n_6_795), .A2 (n_6_1_694));
NAND2_X1 CLOCK_slo__sro_c60698 (.ZN (CLOCK_slo__sro_n55169), .A1 (CLOCK_slo__sro_n55170), .A2 (CLOCK_slo__sro_n55171));
BUF_X4 spw__c75087 (.Z (slo__n5306), .A (spw__n66887));
NAND2_X1 CLOCK_slo__sro_c60681 (.ZN (CLOCK_slo__sro_n55157), .A1 (n_6_1_764), .A2 (n_6_649));
NAND2_X1 CLOCK_slo__sro_c60682 (.ZN (CLOCK_slo__sro_n55156), .A1 (CLOCK_slo__sro_n55157), .A2 (slo__sro_n27862));
AOI21_X2 CLOCK_slo__sro_c60683 (.ZN (slo__sro_n27860), .A (CLOCK_slo__sro_n55156)
    , .B1 (n_6_681), .B2 (n_6_1_765));
INV_X1 CLOCK_slo__c60830 (.ZN (CLOCK_slo__n55287), .A (n_6_1_547));
INV_X2 CLOCK_slo__c60932 (.ZN (CLOCK_slo__n55377), .A (slo__sro_n27836));
INV_X1 CLOCK_slo__sro_c61440 (.ZN (CLOCK_slo__sro_n55809), .A (CLOCK_sgo__n46934));
INV_X1 CLOCK_slo__c61094 (.ZN (CLOCK_slo__n55511), .A (n_6_1_504));
INV_X1 CLOCK_slo__c60766 (.ZN (CLOCK_slo__n55232), .A (n_6_1_825));
INV_X2 CLOCK_slo__c61380 (.ZN (CLOCK_slo__n55755), .A (slo__sro_n34606));
NAND2_X2 CLOCK_slo__sro_c60960 (.ZN (CLOCK_slo__sro_n55399), .A1 (n_6_609), .A2 (n_6_1_800));
INV_X1 CLOCK_slo__c60861 (.ZN (CLOCK_slo__n55312), .A (slo__sro_n17646));
INV_X2 CLOCK_slo__c61242 (.ZN (CLOCK_slo__n55647), .A (n_6_1_792));
NAND2_X1 CLOCK_slo__sro_c60959 (.ZN (CLOCK_slo__sro_n55400), .A1 (n_6_2636), .A2 (n_6_1_798));
NAND2_X2 CLOCK_slo__sro_c60961 (.ZN (CLOCK_slo__sro_n55398), .A1 (CLOCK_slo__sro_n55399), .A2 (CLOCK_slo__sro_n55400));
AOI21_X2 CLOCK_slo__sro_c60962 (.ZN (n_6_1_767), .A (CLOCK_slo__sro_n55398), .B1 (n_6_577), .B2 (n_6_1_799));
NAND2_X1 CLOCK_slo__sro_c61012 (.ZN (CLOCK_slo__sro_n55449), .A1 (n_6_165), .A2 (n_6_1_1045));
AOI21_X1 CLOCK_slo__sro_c61013 (.ZN (CLOCK_slo__sro_n55448), .A (slo__sro_n34247)
    , .B1 (n_6_133), .B2 (n_6_1_1044));
AND2_X2 CLOCK_slo__sro_c61014 (.ZN (CLOCK_slo__sro_n55447), .A1 (CLOCK_slo__sro_n55448), .A2 (CLOCK_slo__sro_n55449));
NOR2_X1 CLOCK_slo__sro_c61441 (.ZN (CLOCK_slo__sro_n55808), .A1 (CLOCK_slo__sro_n55810), .A2 (CLOCK_slo__sro_n55809));
AOI221_X2 CLOCK_slo__sro_c61442 (.ZN (n_6_1_871), .A (CLOCK_slo__sro_n55808), .B1 (n_6_416)
    , .B2 (n_6_1_905), .C1 (n_6_384), .C2 (n_6_1_904));
INV_X1 CLOCK_slo__c61507 (.ZN (CLOCK_slo__n55860), .A (slo__sro_n41830));
INV_X1 CLOCK_slo__c61515 (.ZN (CLOCK_slo__n55865), .A (n_6_1_971));
NAND2_X1 CLOCK_slo__sro_c61542 (.ZN (CLOCK_slo__sro_n55889), .A1 (n_6_227), .A2 (n_6_1_1010));
NAND2_X1 CLOCK_slo__sro_c61543 (.ZN (CLOCK_slo__sro_n55888), .A1 (CLOCK_slo__sro_n55889), .A2 (CLOCK_slo__sro_n55890));
AOI21_X2 CLOCK_slo__sro_c61544 (.ZN (n_6_1_979), .A (CLOCK_slo__sro_n55888), .B1 (n_6_195), .B2 (n_6_1_1009));
INV_X1 CLOCK_slo__sro_c61603 (.ZN (CLOCK_slo__sro_n55929), .A (CLOCK_slo__sro_n55930));
AND2_X1 CLOCK_slo__sro_c61415 (.ZN (CLOCK_slo__sro_n55785), .A1 (n_6_2623), .A2 (n_6_1_763));
AOI221_X2 CLOCK_slo__sro_c61416 (.ZN (CLOCK_slo__sro_n55784), .A (CLOCK_slo__sro_n55785)
    , .B1 (n_6_659), .B2 (n_6_1_764), .C1 (n_6_691), .C2 (n_6_1_765));
AOI221_X2 CLOCK_slo__sro_c61604 (.ZN (n_6_1_806), .A (CLOCK_slo__sro_n55929), .B1 (n_6_549)
    , .B2 (n_6_1_835), .C1 (n_6_517), .C2 (n_6_1_834));
AND2_X1 CLOCK_slo__sro_c61636 (.ZN (CLOCK_slo__sro_n55959), .A1 (n_6_462), .A2 (n_6_1_869));
NAND2_X2 CLOCK_slo__sro_c61592 (.ZN (slo__sro_n27691), .A1 (n_6_730), .A2 (n_6_1_729));
NAND2_X1 CLOCK_slo__sro_c61709 (.ZN (CLOCK_slo__sro_n56018), .A1 (n_6_181), .A2 (n_6_1_1045));
NAND2_X1 CLOCK_slo__sro_c61710 (.ZN (CLOCK_slo__sro_n56017), .A1 (CLOCK_slo__sro_n56019), .A2 (CLOCK_slo__sro_n56018));
AOI21_X1 CLOCK_slo__sro_c61711 (.ZN (n_6_1_1032), .A (CLOCK_slo__sro_n56017), .B1 (n_6_149), .B2 (n_6_1_1044));
NAND2_X2 CLOCK_slo__sro_c61764 (.ZN (CLOCK_slo__sro_n56058), .A1 (CLOCK_slo__sro_n56059), .A2 (CLOCK_slo__sro_n56060));
AOI21_X2 CLOCK_slo__sro_c61765 (.ZN (CLOCK_slo__sro_n56057), .A (CLOCK_slo__sro_n56058)
    , .B1 (n_6_244), .B2 (n_6_1_1010));
INV_X1 CLOCK_slo__c61787 (.ZN (CLOCK_slo__n56075), .A (n_6_1_1103));
INV_X2 CLOCK_slo__c61974 (.ZN (CLOCK_slo__n56237), .A (slo__sro_n27689));
NOR2_X1 CLOCK_slo__sro_c61736 (.ZN (n_6_1_864), .A1 (slo__sro_n29489), .A2 (CLOCK_slo__sro_n56037));
NAND2_X1 CLOCK_slo__sro_c61763 (.ZN (CLOCK_slo__sro_n56059), .A1 (n_6_212), .A2 (n_6_1_1009));
INV_X1 CLOCK_slo__c61966 (.ZN (CLOCK_slo__n56232), .A (slo__sro_n35183));
AOI222_X2 CLOCK_slo__sro_c61850 (.ZN (CLOCK_slo__sro_n56126), .A1 (n_6_548), .A2 (n_6_1_835)
    , .B1 (n_6_516), .B2 (n_6_1_834), .C1 (n_6_2670), .C2 (CLOCK_sgo__n46922));
NAND2_X1 CLOCK_slo__sro_c61997 (.ZN (CLOCK_slo__sro_n56261), .A1 (n_6_2470), .A2 (n_6_1_588));
INV_X1 CLOCK_slo__sro_c61998 (.ZN (CLOCK_slo__sro_n56260), .A (CLOCK_slo__sro_n56261));
AOI221_X2 CLOCK_slo__sro_c61999 (.ZN (n_6_1_577), .A (CLOCK_slo__sro_n56260), .B1 (n_6_1013)
    , .B2 (slo___n23218), .C1 (n_6_981), .C2 (slo___n23232));
NAND2_X1 CLOCK_slo__sro_c62451 (.ZN (CLOCK_slo__sro_n56610), .A1 (n_6_150), .A2 (n_6_1_1044));
INV_X2 CLOCK_slo__c62070 (.ZN (CLOCK_slo__n56313), .A (slo__sro_n11796));
NAND2_X1 CLOCK_slo__sro_c62147 (.ZN (CLOCK_slo__sro_n56377), .A1 (CLOCK_slo__sro_n56378), .A2 (CLOCK_slo__sro_n56379));
AOI21_X1 CLOCK_slo__sro_c62148 (.ZN (CLOCK_slo__sro_n56376), .A (CLOCK_slo__sro_n56377)
    , .B1 (n_6_566), .B2 (n_6_1_835));
NAND2_X1 CLOCK_slo__sro_c62436 (.ZN (CLOCK_slo__sro_n56597), .A1 (n_6_1_834), .A2 (n_6_538));
INV_X2 CLOCK_slo__c62205 (.ZN (CLOCK_slo__n56418), .A (slo__sro_n29857));
NAND2_X1 CLOCK_slo__sro_c62437 (.ZN (CLOCK_slo__sro_n56596), .A1 (CLOCK_slo__sro_n56597), .A2 (CLOCK_slo__sro_n56598));
AOI21_X1 CLOCK_slo__sro_c62438 (.ZN (n_6_1_827), .A (CLOCK_slo__sro_n56596), .B1 (n_6_570), .B2 (n_6_1_835));
AND2_X1 CLOCK_slo__sro_c62453 (.ZN (CLOCK_slo__sro_n56608), .A1 (CLOCK_slo__sro_n56609), .A2 (CLOCK_slo__sro_n56610));
AOI222_X2 CLOCK_slo__sro_c62667 (.ZN (n_6_1_802), .A1 (n_6_545), .A2 (n_6_1_835), .B1 (n_6_513)
    , .B2 (n_6_1_834), .C1 (n_6_2667), .C2 (CLOCK_sgo__n46922));
INV_X2 CLOCK_slo__c62574 (.ZN (CLOCK_slo__n56713), .A (n_6_1_931));
NOR2_X2 CLOCK_slo__sro_c62634 (.ZN (n_6_1_819), .A1 (slo__sro_n8764), .A2 (CLOCK_slo__sro_n56757));
NAND2_X1 CLOCK_slo__sro_c62810 (.ZN (CLOCK_slo__sro_n56894), .A1 (CLOCK_slo__sro_n56895), .A2 (CLOCK_slo__sro_n56896));
AOI21_X1 CLOCK_slo__sro_c62811 (.ZN (n_6_1_180), .A (CLOCK_slo__sro_n56894), .B1 (n_6_1705), .B2 (slo___n23407));
INV_X1 CLOCK_slo__c62279 (.ZN (CLOCK_slo__n56467), .A (slo__sro_n6955));
NAND2_X1 CLOCK_slo__sro_c63139 (.ZN (CLOCK_slo__sro_n57156), .A1 (CLOCK_opt_ipo_n46038), .A2 (CLOCK_sgo__n46922));
INV_X1 CLOCK_slo__c62889 (.ZN (CLOCK_slo__n56953), .A (slo__sro_n8646));
INV_X1 CLOCK_slo__c62879 (.ZN (CLOCK_slo__n56946), .A (n_6_1_719));
INV_X1 CLOCK_slo__c62610 (.ZN (CLOCK_slo__n56734), .A (slo__sro_n35288));
INV_X2 CLOCK_slo__c62792 (.ZN (CLOCK_slo__n56881), .A (n_6_1_1054));
INV_X1 CLOCK_slo__c62863 (.ZN (CLOCK_slo__n56933), .A (n_6_1_682));
NAND2_X1 CLOCK_slo__sro_c63140 (.ZN (CLOCK_slo__sro_n57155), .A1 (n_6_1_835), .A2 (n_6_552));
NAND2_X1 CLOCK_slo__sro_c63141 (.ZN (CLOCK_slo__sro_n57154), .A1 (CLOCK_slo__sro_n57155), .A2 (CLOCK_slo__sro_n57156));
INV_X1 CLOCK_slo__xsl_c62979 (.ZN (CLOCK_slo__xsl_n57029), .A (slo__sro_n41807));
BUF_X2 CLOCK_slo__xsl_c62981 (.Z (slo___n13100), .A (slo__sro_n41807));
AOI222_X2 CLOCK_slo__sro_c63113 (.ZN (CLOCK_slo__sro_n57132), .A1 (n_6_1866), .A2 (CLOCK_sgo__n48011)
    , .B1 (n_6_1898), .B2 (n_6_1_100), .C1 (n_6_2025), .C2 (n_6_1_98));
AOI221_X2 CLOCK_slo__sro_c63527 (.ZN (slo__sro_n31830), .A (slo__sro_n31831), .B1 (n_6_202)
    , .B2 (n_6_1_1009), .C1 (n_6_234), .C2 (n_6_1_1010));
INV_X1 CLOCK_slo__c63551 (.ZN (CLOCK_slo__n57456), .A (n_6_1_946));
AOI222_X2 CLOCK_slo__sro_c63380 (.ZN (n_6_1_187), .A1 (n_6_1712), .A2 (slo___n23407)
    , .B1 (n_6_1680), .B2 (n_6_1_204), .C1 (n_6_2124), .C2 (n_6_1_203));
INV_X2 CLOCK_slo__c63629 (.ZN (CLOCK_slo__n57518), .A (slo__sro_n19076));
INV_X1 CLOCK_slo__c63584 (.ZN (CLOCK_slo__n57483), .A (CLOCK_slo__sro_n62530));
INV_X2 CLOCK_slo__c63637 (.ZN (CLOCK_slo__n57523), .A (n_6_1_945));
INV_X2 CLOCK_slo__c63682 (.ZN (CLOCK_slo__n57556), .A (CLOCK_slo__sro_n53015));
INV_X1 CLOCK_slo__c63651 (.ZN (CLOCK_slo__n57534), .A (n_6_1_1100));
NAND2_X1 CLOCK_slo__sro_c69873 (.ZN (CLOCK_slo__sro_n62930), .A1 (CLOCK_slo__sro_n62931), .A2 (CLOCK_slo__sro_n62932));
INV_X1 CLOCK_slo__sro_c63882 (.ZN (CLOCK_slo__sro_n57702), .A (n_6_1_272));
INV_X2 CLOCK_slo__c63670 (.ZN (CLOCK_slo__n57547), .A (slo__sro_n12865));
NAND2_X1 CLOCK_slo__sro_c63868 (.ZN (CLOCK_slo__sro_n57687), .A1 (CLOCK_opt_ipo_n45969), .A2 (n_6_1_273));
INV_X1 CLOCK_slo__sro_c63869 (.ZN (CLOCK_slo__sro_n57686), .A (CLOCK_slo__sro_n57687));
AOI221_X2 CLOCK_slo__sro_c63870 (.ZN (CLOCK_slo__sro_n57685), .A (CLOCK_slo__sro_n57686)
    , .B1 (n_6_1573), .B2 (slo___n23244), .C1 (n_6_1541), .C2 (n_6_1_274));
BUF_X1 spt__c74617 (.Z (n_6_1_182), .A (spt__n66415));
INV_X2 CLOCK_slo__c64155 (.ZN (CLOCK_slo__n57906), .A (n_6_1_540));
INV_X1 CLOCK_slo__c64015 (.ZN (CLOCK_slo__n57799), .A (n_6_1_439));
INV_X1 CLOCK_slo__c64256 (.ZN (CLOCK_slo__n57977), .A (CLOCK_slo__sro_n61394));
INV_X2 CLOCK_slo__c63967 (.ZN (CLOCK_slo__n57760), .A (CLOCK_sgo__sro_n47835));
INV_X2 CLOCK_slo__c64142 (.ZN (CLOCK_slo__n57899), .A (slo__sro_n28333));
AOI221_X2 CLOCK_slo__sro_c64883 (.ZN (n_6_1_93), .A (CLOCK_slo__sro_n58465), .B1 (n_6_1883)
    , .B2 (CLOCK_sgo__n48011), .C1 (n_6_1915), .C2 (n_6_1_100));
INV_X2 CLOCK_slo__c64411 (.ZN (CLOCK_slo__n58099), .A (slo__sro_n39363));
INV_X2 CLOCK_slo__c64108 (.ZN (CLOCK_slo__n57874), .A (slo__sro_n4774));
INV_X1 CLOCK_slo__sro_c64460 (.ZN (CLOCK_slo__sro_n58146), .A (slo__sro_n34035));
NAND2_X1 CLOCK_slo__sro_c64461 (.ZN (CLOCK_slo__sro_n58145), .A1 (n_6_1_765), .A2 (n_6_687));
NAND2_X1 CLOCK_slo__sro_c64462 (.ZN (CLOCK_slo__sro_n58144), .A1 (CLOCK_slo__sro_n58145), .A2 (CLOCK_slo__sro_n58146));
INV_X2 CLOCK_slo__c63944 (.ZN (CLOCK_slo__n57743), .A (slo__sro_n39249));
AOI21_X2 CLOCK_slo__sro_c64463 (.ZN (slo__sro_n34034), .A (CLOCK_slo__sro_n58144)
    , .B1 (n_6_655), .B2 (n_6_1_764));
NAND2_X1 CLOCK_slo__sro_c64710 (.ZN (CLOCK_slo__sro_n58342), .A1 (n_6_264), .A2 (n_6_1_974));
INV_X2 CLOCK_slo__c64527 (.ZN (CLOCK_slo__n58195), .A (CLOCK_slo__sro_n49672));
AOI221_X2 CLOCK_slo__sro_c64597 (.ZN (n_6_1_88), .A (CLOCK_slo__sro_n49937), .B1 (n_6_1910)
    , .B2 (n_6_1_100), .C1 (n_6_1878), .C2 (CLOCK_sgo__n48011));
AOI21_X1 CLOCK_slo__sro_c64712 (.ZN (n_6_1_949), .A (CLOCK_slo__sro_n58341), .B1 (n_6_296), .B2 (n_6_1_975));
NAND2_X1 CLOCK_slo__sro_c64566 (.ZN (CLOCK_slo__sro_n58235), .A1 (n_6_1_308), .A2 (n_6_2202));
INV_X1 CLOCK_slo__sro_c64567 (.ZN (CLOCK_slo__sro_n58234), .A (CLOCK_slo__sro_n58235));
AOI221_X2 CLOCK_slo__sro_c64568 (.ZN (slo__sro_n36260), .A (CLOCK_slo__sro_n58234)
    , .B1 (n_6_1505), .B2 (slo___n23247), .C1 (n_6_1473), .C2 (n_6_1_309));
INV_X1 CLOCK_slo__sro_c64676 (.ZN (CLOCK_slo__sro_n58314), .A (CLOCK_slo__sro_n58315));
AOI221_X2 CLOCK_slo__sro_c64677 (.ZN (CLOCK_slo__sro_n58313), .A (CLOCK_slo__sro_n58314)
    , .B1 (n_6_611), .B2 (n_6_1_800), .C1 (n_6_579), .C2 (n_6_1_799));
CLKBUF_X1 CLOCK_slo___L1_c1_c64786 (.Z (n_6_2759), .A (CLOCK_slo___n58400));
INV_X1 CLOCK_slo__c64820 (.ZN (CLOCK_slo__n58422), .A (n_6_1_1029));
NAND2_X1 CLOCK_slo__sro_c65145 (.ZN (CLOCK_slo__sro_n58699), .A1 (n_6_610), .A2 (n_6_1_800));
NAND2_X1 CLOCK_slo__sro_c65050 (.ZN (CLOCK_slo__sro_n58611), .A1 (n_6_1_378), .A2 (CLOCK_opt_ipo_n45906));
CLKBUF_X2 spw__c75002 (.Z (slo__sro_n36849), .A (spw__n66802));
AND2_X2 CLOCK_slo__sro_c69434 (.ZN (CLOCK_slo__sro_n62531), .A1 (n_6_80), .A2 (n_6_1_1079));
NAND2_X1 CLOCK_slo__sro_c65146 (.ZN (CLOCK_slo__sro_n58698), .A1 (CLOCK_slo__sro_n58699), .A2 (CLOCK_slo__sro_n58700));
AOI21_X2 CLOCK_slo__sro_c65147 (.ZN (slo__sro_n40959), .A (CLOCK_slo__sro_n58698)
    , .B1 (n_6_578), .B2 (n_6_1_799));
AOI21_X2 CLOCK_slo__sro_c65161 (.ZN (CLOCK_slo__sro_n58708), .A (CLOCK_slo__sro_n58709)
    , .B1 (n_6_1658), .B2 (drc_ipo_n26601));
NAND2_X1 CLOCK_slo__sro_c65216 (.ZN (CLOCK_slo__sro_n58765), .A1 (n_6_1171), .A2 (slo___n23364));
NAND2_X1 CLOCK_slo__sro_c65217 (.ZN (CLOCK_slo__sro_n58764), .A1 (CLOCK_slo__sro_n58765), .A2 (CLOCK_slo__sro_n58766));
AOI21_X2 CLOCK_slo__sro_c65218 (.ZN (n_6_1_470), .A (CLOCK_slo__sro_n58764), .B1 (n_6_1203), .B2 (slo___n23466));
NAND2_X1 CLOCK_slo__sro_c65307 (.ZN (CLOCK_slo__sro_n58847), .A1 (n_6_916), .A2 (slo___n23367));
INV_X1 CLOCK_slo__sro_c64948 (.ZN (CLOCK_slo__sro_n58521), .A (slo__sro_n7436));
AND2_X1 CLOCK_slo__sro_c64949 (.ZN (CLOCK_slo__sro_n58520), .A1 (n_6_1127), .A2 (slo___n23268));
NAND2_X1 CLOCK_slo__sro_c64950 (.ZN (CLOCK_slo__sro_n58519), .A1 (n_6_1095), .A2 (slo___n23277));
NAND2_X1 CLOCK_slo__sro_c64951 (.ZN (CLOCK_slo__sro_n58518), .A1 (CLOCK_slo__sro_n58519), .A2 (CLOCK_slo__sro_n58521));
NOR2_X2 CLOCK_slo__sro_c64952 (.ZN (slo__sro_n7435), .A1 (CLOCK_slo__sro_n58520), .A2 (CLOCK_slo__sro_n58518));
AOI21_X2 CLOCK_slo__sro_c65309 (.ZN (n_6_1_611), .A (CLOCK_slo__sro_n58846), .B1 (n_6_948), .B2 (n_6_1_625));
INV_X1 CLOCK_slo__sro_c65371 (.ZN (CLOCK_slo__sro_n58907), .A (slo__sro_n17598));
NAND2_X1 CLOCK_slo__sro_c65372 (.ZN (CLOCK_slo__sro_n58906), .A1 (n_6_1114), .A2 (slo___n23277));
NAND2_X1 CLOCK_slo__sro_c65373 (.ZN (CLOCK_slo__sro_n58905), .A1 (CLOCK_slo__sro_n58906), .A2 (CLOCK_slo__sro_n58907));
AOI21_X2 CLOCK_slo__sro_c65374 (.ZN (CLOCK_slo__sro_n58904), .A (CLOCK_slo__sro_n58905)
    , .B1 (n_6_1146), .B2 (slo___n23268));
NAND2_X1 CLOCK_slo__sro_c65774 (.ZN (CLOCK_slo__sro_n59282), .A1 (n_6_238), .A2 (n_6_1_1010));
NAND2_X1 CLOCK_slo__sro_c65775 (.ZN (CLOCK_slo__sro_n59281), .A1 (CLOCK_slo__sro_n59282), .A2 (CLOCK_slo__sro_n59283));
INV_X1 CLOCK_slo__sro_c65529 (.ZN (CLOCK_slo__sro_n59058), .A (slo__sro_n9948));
NAND2_X1 CLOCK_slo__sro_c65530 (.ZN (CLOCK_slo__sro_n59057), .A1 (n_6_667), .A2 (n_6_1_764));
NAND2_X1 CLOCK_slo__sro_c65531 (.ZN (CLOCK_slo__sro_n59056), .A1 (CLOCK_slo__sro_n59057), .A2 (CLOCK_slo__sro_n59058));
AOI21_X2 CLOCK_slo__sro_c65532 (.ZN (slo__n35733), .A (CLOCK_slo__sro_n59056), .B1 (n_6_699), .B2 (n_6_1_765));
NAND2_X1 CLOCK_slo__sro_c65608 (.ZN (CLOCK_slo__sro_n59128), .A1 (n_6_1_869), .A2 (n_6_456));
NAND2_X1 CLOCK_slo__sro_c65609 (.ZN (CLOCK_slo__sro_n59127), .A1 (CLOCK_slo__sro_n59128), .A2 (CLOCK_sgo__sro_n47307));
AOI21_X2 CLOCK_slo__sro_c65610 (.ZN (CLOCK_slo__sro_n59126), .A (CLOCK_slo__sro_n59127)
    , .B1 (n_6_488), .B2 (n_6_1_870));
INV_X1 CLOCK_slo__sro_c65796 (.ZN (CLOCK_slo__sro_n59303), .A (CLOCK_slo__sro_n59304));
CLKBUF_X1 spw__L2_c2_c77589 (.Z (n_6_2097), .A (spw__n69100));
AND2_X1 CLOCK_slo__sro_c69952 (.ZN (CLOCK_slo__sro_n63005), .A1 (n_6_2435), .A2 (n_6_1_553));
NAND2_X1 CLOCK_slo__sro_c65501 (.ZN (CLOCK_slo__sro_n59029), .A1 (n_6_305), .A2 (n_6_1_975));
NAND2_X1 CLOCK_slo__sro_c65502 (.ZN (CLOCK_slo__sro_n59028), .A1 (slo__sro_n21836), .A2 (CLOCK_slo__sro_n59029));
AOI21_X2 CLOCK_slo__sro_c65503 (.ZN (CLOCK_slo__sro_n59027), .A (CLOCK_slo__sro_n59028)
    , .B1 (n_6_273), .B2 (n_6_1_974));
NAND2_X1 CLOCK_slo__sro_c65840 (.ZN (CLOCK_slo__sro_n59343), .A1 (CLOCK_slo__sro_n59344), .A2 (CLOCK_slo__sro_n59345));
AOI21_X2 CLOCK_slo__sro_c65841 (.ZN (CLOCK_slo__sro_n59342), .A (CLOCK_slo__sro_n59343)
    , .B1 (n_6_914), .B2 (slo___n23367));
AOI221_X2 CLOCK_slo__sro_c65943 (.ZN (n_6_1_335), .A (CLOCK_slo__sro_n59437), .B1 (n_6_1432)
    , .B2 (slo___n23229), .C1 (n_6_1464), .C2 (n_6_1_345));
AOI221_X2 CLOCK_slo__sro_c65957 (.ZN (CLOCK_slo__sro_n59447), .A (CLOCK_slo__sro_n59448)
    , .B1 (n_6_1494), .B2 (n_6_1_309), .C1 (n_6_1526), .C2 (slo___n23247));
NAND2_X1 CLOCK_slo__sro_c65979 (.ZN (CLOCK_slo__sro_n59469), .A1 (slo__n30670), .A2 (n_6_1_483));
NAND2_X1 CLOCK_slo__sro_c65980 (.ZN (CLOCK_slo__sro_n59468), .A1 (n_6_1159), .A2 (slo___n23364));
NAND2_X1 CLOCK_slo__sro_c65981 (.ZN (CLOCK_slo__sro_n59467), .A1 (CLOCK_slo__sro_n59468), .A2 (CLOCK_slo__sro_n59469));
AOI21_X2 CLOCK_slo__sro_c65982 (.ZN (n_6_1_458), .A (CLOCK_slo__sro_n59467), .B1 (n_6_1191), .B2 (slo___n23466));
NAND2_X1 CLOCK_slo__sro_c66054 (.ZN (CLOCK_slo__sro_n59533), .A1 (CLOCK_slo__sro_n59534), .A2 (CLOCK_slo__sro_n59535));
AOI21_X2 CLOCK_slo__sro_c66055 (.ZN (slo__sro_n13278), .A (CLOCK_slo__sro_n59533)
    , .B1 (n_6_1745), .B2 (n_6_1_169));
INV_X1 CLOCK_slo__sro_c66073 (.ZN (CLOCK_slo__sro_n59550), .A (CLOCK_slo__sro_n59551));
AOI221_X1 CLOCK_slo__sro_c66074 (.ZN (CLOCK_slo__sro_n59549), .A (CLOCK_slo__sro_n59550)
    , .B1 (n_6_1409), .B2 (slo___n23229), .C1 (n_6_1441), .C2 (n_6_1_345));
NOR2_X2 CLOCK_slo__sro_c66168 (.ZN (slo__sro_n6762), .A1 (slo__sro_n6763), .A2 (CLOCK_slo__sro_n59641));
NAND2_X1 CLOCK_slo__sro_c66246 (.ZN (CLOCK_slo__sro_n59714), .A1 (n_6_2787), .A2 (CLOCK_sgo__n46937));
INV_X1 CLOCK_slo__sro_c66247 (.ZN (CLOCK_slo__sro_n59713), .A (CLOCK_slo__sro_n59714));
AOI221_X2 CLOCK_slo__sro_c66248 (.ZN (CLOCK_slo__sro_n59712), .A (CLOCK_slo__sro_n59713)
    , .B1 (n_6_348), .B2 (n_6_1_939), .C1 (n_6_380), .C2 (n_6_1_940));
NAND2_X1 CLOCK_slo__sro_c66264 (.ZN (CLOCK_slo__sro_n59728), .A1 (CLOCK_slo__sro_n59729), .A2 (CLOCK_slo__sro_n59730));
AOI21_X2 CLOCK_slo__sro_c66265 (.ZN (slo__sro_n39249), .A (CLOCK_slo__sro_n59728)
    , .B1 (n_6_1879), .B2 (CLOCK_sgo__n48011));
NOR2_X2 CLOCK_slo__sro_c66506 (.ZN (slo__sro_n12923), .A1 (CLOCK_slo__sro_n59951), .A2 (slo__sro_n12924));
AOI21_X1 CLOCK_slo__sro_c66520 (.ZN (CLOCK_slo__sro_n59961), .A (slo__sro_n22432)
    , .B1 (n_6_272), .B2 (n_6_1_974));
AND2_X1 CLOCK_slo__sro_c66521 (.ZN (slo__sro_n22431), .A1 (CLOCK_slo__sro_n59961), .A2 (CLOCK_slo__sro_n59962));
INV_X1 CLOCK_slo__sro_c66622 (.ZN (CLOCK_slo__sro_n60053), .A (CLOCK_slo__sro_n60054));
NAND2_X1 CLOCK_slo__sro_c66384 (.ZN (CLOCK_slo__sro_n59845), .A1 (n_6_2518), .A2 (n_6_1_658));
NAND2_X1 CLOCK_slo__sro_c66385 (.ZN (CLOCK_slo__sro_n59844), .A1 (n_6_839), .A2 (slo___n23463));
NAND2_X1 CLOCK_slo__sro_c66386 (.ZN (CLOCK_slo__sro_n59843), .A1 (CLOCK_slo__sro_n59844), .A2 (CLOCK_slo__sro_n59845));
NAND2_X1 CLOCK_slo__sro_c66314 (.ZN (CLOCK_slo__sro_n59775), .A1 (n_6_335), .A2 (n_6_1_939));
AOI21_X1 CLOCK_slo__sro_c66315 (.ZN (CLOCK_slo__sro_n59774), .A (slo__sro_n5353), .B1 (n_6_367), .B2 (n_6_1_940));
AND2_X1 CLOCK_slo__sro_c66316 (.ZN (CLOCK_slo__sro_n59773), .A1 (CLOCK_slo__sro_n59774), .A2 (CLOCK_slo__sro_n59775));
INV_X1 CLOCK_slo__sro_c66705 (.ZN (CLOCK_slo__sro_n60126), .A (CLOCK_slo__sro_n60127));
NOR2_X1 CLOCK_slo__sro_c66706 (.ZN (CLOCK_slo__sro_n60125), .A1 (slo__sro_n37306), .A2 (CLOCK_slo__sro_n60126));
NAND2_X1 CLOCK_slo__sro_c66878 (.ZN (CLOCK_slo__sro_n60277), .A1 (n_6_1_835), .A2 (n_6_560));
NAND2_X1 CLOCK_slo__sro_c66879 (.ZN (CLOCK_slo__sro_n60276), .A1 (CLOCK_slo__sro_n60277), .A2 (CLOCK_slo__sro_n60278));
AOI21_X1 CLOCK_slo__sro_c66880 (.ZN (CLOCK_slo__sro_n60275), .A (CLOCK_slo__sro_n60276)
    , .B1 (n_6_528), .B2 (n_6_1_834));
INV_X8 CLOCK_slo__c67284 (.ZN (CLOCK_slo__n60587), .A (CLOCK_slo__n60586));
AND2_X2 CLOCK_slo__sro_c66917 (.ZN (CLOCK_slo__sro_n60310), .A1 (n_6_1722), .A2 (slo___n23407));
NOR2_X4 CLOCK_slo__sro_c66918 (.ZN (CLOCK_slo__sro_n60309), .A1 (slo__sro_n38941), .A2 (CLOCK_slo__sro_n60310));
NAND2_X1 CLOCK_slo__sro_c67302 (.ZN (CLOCK_slo__sro_n60605), .A1 (n_6_1833), .A2 (n_6_1_135));
NAND2_X1 CLOCK_slo__sro_c67303 (.ZN (CLOCK_slo__sro_n60604), .A1 (slo__sro_n10694), .A2 (CLOCK_slo__sro_n60605));
AOI21_X2 CLOCK_slo__sro_c67304 (.ZN (CLOCK_slo__sro_n60603), .A (CLOCK_slo__sro_n60604)
    , .B1 (n_6_1801), .B2 (n_6_1_134));
NAND2_X1 CLOCK_slo__sro_c67393 (.ZN (CLOCK_slo__sro_n60681), .A1 (n_6_378), .A2 (n_6_1_940));
INV_X1 CLOCK_slo__sro_c67340 (.ZN (CLOCK_slo__sro_n60642), .A (n_6_1974));
INV_X1 CLOCK_slo__sro_c67341 (.ZN (CLOCK_slo__sro_n60641), .A (n_6_1_65));
NAND2_X1 CLOCK_slo__sro_c67342 (.ZN (CLOCK_slo__sro_n60640), .A1 (n_6_2006), .A2 (n_6_1_63));
OAI21_X1 CLOCK_slo__sro_c67343 (.ZN (CLOCK_slo__sro_n60639), .A (CLOCK_slo__sro_n60640)
    , .B1 (CLOCK_slo__sro_n60642), .B2 (CLOCK_slo__sro_n60641));
AOI21_X1 CLOCK_slo__sro_c67344 (.ZN (n_6_1_53), .A (CLOCK_slo__sro_n60639), .B1 (n_6_1942), .B2 (n_6_1_64));
AND2_X1 CLOCK_slo__sro_c67395 (.ZN (CLOCK_slo__sro_n60679), .A1 (CLOCK_slo__sro_n60681), .A2 (CLOCK_slo__sro_n60680));
NAND2_X1 CLOCK_slo__sro_c67498 (.ZN (CLOCK_slo__sro_n60777), .A1 (n_6_1735), .A2 (n_6_1_169));
NAND2_X1 CLOCK_slo__sro_c67499 (.ZN (CLOCK_slo__sro_n60776), .A1 (CLOCK_slo__sro_n60777), .A2 (CLOCK_slo__sro_n60778));
AOI21_X2 CLOCK_slo__sro_c67500 (.ZN (n_6_1_143), .A (CLOCK_slo__sro_n60776), .B1 (n_6_1767), .B2 (n_6_1_170));
NAND2_X1 CLOCK_slo__sro_c67542 (.ZN (CLOCK_slo__sro_n60814), .A1 (n_6_1681), .A2 (n_6_1_204));
NAND2_X1 CLOCK_slo__sro_c67543 (.ZN (CLOCK_slo__sro_n60813), .A1 (n_6_1713), .A2 (slo___n23407));
AND3_X1 CLOCK_slo__sro_c67544 (.ZN (CLOCK_slo__sro_n60812), .A1 (CLOCK_slo__sro_n60814)
    , .A2 (CLOCK_slo__sro_n60815), .A3 (CLOCK_slo__sro_n60813));
INV_X4 CLOCK_slo__c67583 (.ZN (slo__sro_n14967), .A (CLOCK_slo__n60839));

endmodule //BoothAlgorithmMultiplier

module BAMIntegrated (clk, Multiplicand, Multiplier, enableA, enableB, enableOut, 
    resetA, resetB, resetOut, Product);

output [63:0] Product;
input [31:0] Multiplicand;
input [31:0] Multiplier;
input clk;
input enableA;
input enableB;
input enableOut;
input resetA;
input resetB;
input resetOut;
wire CTS_n618;
wire CLOCK_slh_n790;
wire CLOCK_slh_n800;
wire CLOCK_slh_n845;
wire sph__n1141;
wire sph__n1144;
wire sph__n1163;
wire sph__n1198;
wire sph__n1189;
wire sph__n1201;
wire sph__n1195;
wire sph__n1192;
wire sph__n1207;
wire sph__n1204;
wire CLOCK_slh_n928;
wire sph__n1166;
wire sph__n1169;
wire sph__n1183;
wire sph__n1172;
wire sph__n1186;
wire CLOCK_slh_n840;
wire CLOCK_slh_n870;
wire \registerInProduct[63] ;
wire \registerInProduct[62] ;
wire \registerInProduct[61] ;
wire \registerInProduct[60] ;
wire \registerInProduct[59] ;
wire \registerInProduct[58] ;
wire \registerInProduct[57] ;
wire \registerInProduct[56] ;
wire \registerInProduct[55] ;
wire \registerInProduct[54] ;
wire \registerInProduct[53] ;
wire \registerInProduct[52] ;
wire \registerInProduct[51] ;
wire \registerInProduct[50] ;
wire \registerInProduct[49] ;
wire \registerInProduct[48] ;
wire \registerInProduct[47] ;
wire \registerInProduct[46] ;
wire \registerInProduct[45] ;
wire \registerInProduct[44] ;
wire \registerInProduct[43] ;
wire \registerInProduct[42] ;
wire \registerInProduct[41] ;
wire \registerInProduct[40] ;
wire \registerInProduct[39] ;
wire \registerInProduct[38] ;
wire \registerInProduct[37] ;
wire \registerInProduct[36] ;
wire \registerInProduct[35] ;
wire \registerInProduct[34] ;
wire \registerInProduct[33] ;
wire \registerInProduct[32] ;
wire \registerInProduct[31] ;
wire \registerInProduct[30] ;
wire \registerInProduct[29] ;
wire \registerInProduct[28] ;
wire \registerInProduct[27] ;
wire \registerInProduct[26] ;
wire \registerInProduct[25] ;
wire \registerInProduct[24] ;
wire \registerInProduct[23] ;
wire \registerInProduct[22] ;
wire \registerInProduct[21] ;
wire \registerInProduct[20] ;
wire \registerInProduct[19] ;
wire \registerInProduct[18] ;
wire \registerInProduct[17] ;
wire \registerInProduct[16] ;
wire \registerInProduct[15] ;
wire \registerInProduct[14] ;
wire \registerInProduct[13] ;
wire \registerInProduct[12] ;
wire \registerInProduct[11] ;
wire \registerInProduct[10] ;
wire \registerInProduct[9] ;
wire \registerInProduct[8] ;
wire \registerInProduct[7] ;
wire \registerInProduct[6] ;
wire \registerInProduct[5] ;
wire \registerInProduct[4] ;
wire \registerInProduct[3] ;
wire \registerInProduct[2] ;
wire \registerInProduct[1] ;
wire \registerInProduct[0] ;
wire CTS_n564;
wire \InputRegisterA_register[31] ;
wire \InputRegisterA_register[30] ;
wire \InputRegisterA_register[29] ;
wire \InputRegisterA_register[28] ;
wire \InputRegisterA_register[27] ;
wire \InputRegisterA_register[26] ;
wire \InputRegisterA_register[25] ;
wire \InputRegisterA_register[24] ;
wire \InputRegisterA_register[23] ;
wire \InputRegisterA_register[22] ;
wire \InputRegisterA_register[21] ;
wire \InputRegisterA_register[20] ;
wire \InputRegisterA_register[19] ;
wire \InputRegisterA_register[18] ;
wire \InputRegisterA_register[17] ;
wire \InputRegisterA_register[16] ;
wire \InputRegisterA_register[15] ;
wire \InputRegisterA_register[14] ;
wire \InputRegisterA_register[13] ;
wire \InputRegisterA_register[12] ;
wire \InputRegisterA_register[11] ;
wire \InputRegisterA_register[10] ;
wire \InputRegisterA_register[9] ;
wire \InputRegisterA_register[8] ;
wire \InputRegisterA_register[7] ;
wire \InputRegisterA_register[6] ;
wire \InputRegisterA_register[5] ;
wire \InputRegisterA_register[4] ;
wire \InputRegisterA_register[3] ;
wire \InputRegisterA_register[2] ;
wire \InputRegisterA_register[1] ;
wire \InputRegisterA_register[0] ;
wire \registerOutA[31] ;
wire \registerOutA[30] ;
wire \registerOutA[29] ;
wire \registerOutA[28] ;
wire \registerOutA[27] ;
wire \registerOutA[26] ;
wire \registerOutA[25] ;
wire \registerOutA[24] ;
wire \registerOutA[23] ;
wire \registerOutA[22] ;
wire \registerOutA[21] ;
wire \registerOutA[20] ;
wire \registerOutA[19] ;
wire \registerOutA[18] ;
wire \registerOutA[17] ;
wire \registerOutA[16] ;
wire \registerOutA[15] ;
wire \registerOutA[14] ;
wire \registerOutA[13] ;
wire \registerOutA[12] ;
wire \registerOutA[11] ;
wire \registerOutA[10] ;
wire \registerOutA[9] ;
wire \registerOutA[8] ;
wire \registerOutA[7] ;
wire \registerOutA[6] ;
wire \registerOutA[5] ;
wire \registerOutA[4] ;
wire \registerOutA[3] ;
wire \registerOutA[2] ;
wire drc_ipo_n350;
wire CTS_n560;
wire \InputRegisterB_register[31] ;
wire \InputRegisterB_register[30] ;
wire \InputRegisterB_register[29] ;
wire \InputRegisterB_register[28] ;
wire \InputRegisterB_register[27] ;
wire \InputRegisterB_register[26] ;
wire \InputRegisterB_register[25] ;
wire \InputRegisterB_register[24] ;
wire \InputRegisterB_register[23] ;
wire \InputRegisterB_register[22] ;
wire \InputRegisterB_register[21] ;
wire \InputRegisterB_register[20] ;
wire \InputRegisterB_register[19] ;
wire \InputRegisterB_register[18] ;
wire \InputRegisterB_register[17] ;
wire \InputRegisterB_register[16] ;
wire \InputRegisterB_register[15] ;
wire \InputRegisterB_register[14] ;
wire \InputRegisterB_register[13] ;
wire \InputRegisterB_register[12] ;
wire \InputRegisterB_register[11] ;
wire \InputRegisterB_register[10] ;
wire \InputRegisterB_register[9] ;
wire \InputRegisterB_register[8] ;
wire \InputRegisterB_register[7] ;
wire \InputRegisterB_register[6] ;
wire \InputRegisterB_register[5] ;
wire \InputRegisterB_register[4] ;
wire \InputRegisterB_register[3] ;
wire \InputRegisterB_register[2] ;
wire \InputRegisterB_register[1] ;
wire \InputRegisterB_register[0] ;
wire \registerOutB[31] ;
wire \registerOutB[30] ;
wire \registerOutB[29] ;
wire \registerOutB[28] ;
wire \registerOutB[27] ;
wire \registerOutB[26] ;
wire \registerOutB[25] ;
wire \registerOutB[24] ;
wire \registerOutB[23] ;
wire \registerOutB[22] ;
wire \registerOutB[21] ;
wire \registerOutB[20] ;
wire \registerOutB[19] ;
wire \registerOutB[18] ;
wire \registerOutB[17] ;
wire \registerOutB[16] ;
wire \registerOutB[15] ;
wire \registerOutB[14] ;
wire \registerOutB[13] ;
wire \registerOutB[12] ;
wire \registerOutB[11] ;
wire \registerOutB[10] ;
wire \registerOutB[9] ;
wire \registerOutB[8] ;
wire \registerOutB[7] ;
wire \registerOutB[6] ;
wire \registerOutB[5] ;
wire \registerOutB[4] ;
wire \registerOutB[3] ;
wire \registerOutB[2] ;
wire \registerOutB[1] ;
wire drc_ipo_n348;
wire \OutputRegister_register[63] ;
wire \OutputRegister_register[62] ;
wire \OutputRegister_register[61] ;
wire \OutputRegister_register[60] ;
wire \OutputRegister_register[59] ;
wire \OutputRegister_register[58] ;
wire \OutputRegister_register[57] ;
wire \OutputRegister_register[56] ;
wire \OutputRegister_register[55] ;
wire \OutputRegister_register[54] ;
wire \OutputRegister_register[53] ;
wire \OutputRegister_register[52] ;
wire \OutputRegister_register[51] ;
wire \OutputRegister_register[50] ;
wire \OutputRegister_register[49] ;
wire \OutputRegister_register[48] ;
wire \OutputRegister_register[47] ;
wire \OutputRegister_register[46] ;
wire \OutputRegister_register[45] ;
wire \OutputRegister_register[44] ;
wire \OutputRegister_register[43] ;
wire \OutputRegister_register[42] ;
wire \OutputRegister_register[41] ;
wire \OutputRegister_register[40] ;
wire \OutputRegister_register[39] ;
wire \OutputRegister_register[38] ;
wire \OutputRegister_register[37] ;
wire \OutputRegister_register[36] ;
wire \OutputRegister_register[35] ;
wire \OutputRegister_register[34] ;
wire \OutputRegister_register[33] ;
wire \OutputRegister_register[32] ;
wire \OutputRegister_register[31] ;
wire \OutputRegister_register[30] ;
wire \OutputRegister_register[29] ;
wire \OutputRegister_register[28] ;
wire \OutputRegister_register[27] ;
wire \OutputRegister_register[26] ;
wire \OutputRegister_register[25] ;
wire \OutputRegister_register[24] ;
wire \OutputRegister_register[23] ;
wire \OutputRegister_register[22] ;
wire \OutputRegister_register[21] ;
wire \OutputRegister_register[20] ;
wire \OutputRegister_register[19] ;
wire \OutputRegister_register[18] ;
wire \OutputRegister_register[17] ;
wire \OutputRegister_register[16] ;
wire \OutputRegister_register[15] ;
wire \OutputRegister_register[14] ;
wire \OutputRegister_register[13] ;
wire \OutputRegister_register[12] ;
wire \OutputRegister_register[11] ;
wire \OutputRegister_register[10] ;
wire \OutputRegister_register[9] ;
wire \OutputRegister_register[8] ;
wire \OutputRegister_register[7] ;
wire \OutputRegister_register[6] ;
wire \OutputRegister_register[5] ;
wire \OutputRegister_register[4] ;
wire \OutputRegister_register[3] ;
wire \OutputRegister_register[2] ;
wire \OutputRegister_register[1] ;
wire \OutputRegister_register[0] ;
wire InputRegisterA_n_1;
wire InputRegisterB_n_1;
wire OutputRegister_n_1;
wire CTS_n617;
wire InputRegisterB_n_2;
wire InputRegisterB_n_4;
wire InputRegisterB_n_5;
wire InputRegisterB_n_6;
wire InputRegisterB_n_7;
wire InputRegisterB_n_8;
wire InputRegisterB_n_9;
wire InputRegisterB_n_10;
wire InputRegisterB_n_11;
wire InputRegisterB_n_12;
wire InputRegisterB_n_13;
wire InputRegisterB_n_14;
wire InputRegisterB_n_15;
wire InputRegisterB_n_16;
wire InputRegisterB_n_17;
wire InputRegisterB_n_18;
wire InputRegisterB_n_19;
wire InputRegisterB_n_20;
wire InputRegisterB_n_21;
wire InputRegisterB_n_22;
wire InputRegisterB_n_23;
wire InputRegisterB_n_24;
wire InputRegisterB_n_25;
wire InputRegisterB_n_26;
wire InputRegisterB_n_27;
wire InputRegisterB_n_28;
wire InputRegisterB_n_29;
wire InputRegisterB_n_30;
wire InputRegisterB_n_31;
wire InputRegisterB_n_32;
wire InputRegisterB_n_33;
wire InputRegisterB_n_34;
wire InputRegisterA_n_2;
wire InputRegisterA_n_4;
wire InputRegisterA_n_5;
wire InputRegisterA_n_6;
wire InputRegisterA_n_7;
wire InputRegisterA_n_8;
wire InputRegisterA_n_9;
wire InputRegisterA_n_10;
wire InputRegisterA_n_11;
wire InputRegisterA_n_12;
wire InputRegisterA_n_13;
wire InputRegisterA_n_14;
wire InputRegisterA_n_15;
wire InputRegisterA_n_16;
wire InputRegisterA_n_17;
wire InputRegisterA_n_18;
wire InputRegisterA_n_19;
wire InputRegisterA_n_20;
wire InputRegisterA_n_21;
wire InputRegisterA_n_22;
wire InputRegisterA_n_23;
wire InputRegisterA_n_24;
wire InputRegisterA_n_25;
wire InputRegisterA_n_26;
wire InputRegisterA_n_27;
wire InputRegisterA_n_28;
wire InputRegisterA_n_29;
wire InputRegisterA_n_30;
wire InputRegisterA_n_31;
wire InputRegisterA_n_32;
wire InputRegisterA_n_33;
wire InputRegisterA_n_34;
wire OutputRegister_n_2;
wire OutputRegister_n_4;
wire OutputRegister_n_5;
wire OutputRegister_n_6;
wire OutputRegister_n_7;
wire OutputRegister_n_8;
wire OutputRegister_n_9;
wire OutputRegister_n_10;
wire OutputRegister_n_11;
wire OutputRegister_n_12;
wire OutputRegister_n_13;
wire OutputRegister_n_14;
wire OutputRegister_n_15;
wire OutputRegister_n_16;
wire OutputRegister_n_17;
wire OutputRegister_n_18;
wire OutputRegister_n_19;
wire OutputRegister_n_20;
wire OutputRegister_n_21;
wire OutputRegister_n_22;
wire OutputRegister_n_23;
wire OutputRegister_n_24;
wire OutputRegister_n_25;
wire OutputRegister_n_26;
wire OutputRegister_n_27;
wire OutputRegister_n_28;
wire OutputRegister_n_29;
wire OutputRegister_n_30;
wire OutputRegister_n_31;
wire OutputRegister_n_32;
wire OutputRegister_n_33;
wire OutputRegister_n_34;
wire OutputRegister_n_35;
wire OutputRegister_n_36;
wire OutputRegister_n_37;
wire OutputRegister_n_38;
wire OutputRegister_n_39;
wire OutputRegister_n_40;
wire OutputRegister_n_41;
wire OutputRegister_n_42;
wire OutputRegister_n_43;
wire OutputRegister_n_44;
wire OutputRegister_n_45;
wire OutputRegister_n_46;
wire OutputRegister_n_47;
wire OutputRegister_n_48;
wire OutputRegister_n_49;
wire OutputRegister_n_50;
wire OutputRegister_n_51;
wire OutputRegister_n_52;
wire OutputRegister_n_53;
wire OutputRegister_n_54;
wire OutputRegister_n_55;
wire OutputRegister_n_56;
wire OutputRegister_n_57;
wire OutputRegister_n_58;
wire OutputRegister_n_59;
wire OutputRegister_n_60;
wire OutputRegister_n_61;
wire OutputRegister_n_62;
wire OutputRegister_n_63;
wire OutputRegister_n_64;
wire OutputRegister_n_65;
wire OutputRegister_n_66;
wire hfn_ipo_n71;
wire hfn_ipo_n72;
wire drc_ipo_n347;
wire hfn_ipo_n74;
wire drc_ipo_n105;
wire drc_ipo_n104;
wire drc_ipo_n103;
wire drc_ipo_n102;
wire drc_ipo_n101;
wire drc_ipo_n100;
wire drc_ipo_n99;
wire drc_ipo_n98;
wire drc_ipo_n97;
wire drc_ipo_n96;
wire drc_ipo_n95;
wire drc_ipo_n94;
wire drc_ipo_n93;
wire drc_ipo_n92;
wire drc_ipo_n91;
wire drc_ipo_n90;
wire drc_ipo_n89;
wire drc_ipo_n88;
wire drc_ipo_n87;
wire drc_ipo_n86;
wire drc_ipo_n85;
wire drc_ipo_n84;
wire drc_ipo_n83;
wire drc_ipo_n82;
wire drc_ipo_n80;
wire drc_ipo_n79;
wire drc_ipo_n78;
wire drc_ipo_n351;
wire drc_ipo_n76;
wire drc_ipo_n353;
wire drc_ipo_n354;
wire CTS_n633;
wire sph_n1140;
wire opt_ipo_n299;
wire drc_ipo_n352;
wire CTS_n565;
wire slo___n231;
wire slo__n236;
wire drc_ipo_n355;
wire CTS_n634;
wire CTS_n630;
wire CTS_n631;
wire slo__n198;
wire CTS_n602;
wire CTS_n619;
wire CTS_n603;
wire CTS_n707;
wire sph_n1154;
wire sph_n1162;
wire sph_n1182;
wire sph_n1217;
wire CLOCK_slh__n943;
wire CLOCK_spc__n1018;


MUX2_X1 i_0_1_95 (.Z (OutputRegister_n_66), .A (Product[0]), .B (\OutputRegister_register[0] ), .S (hfn_ipo_n72));
MUX2_X1 i_0_1_94 (.Z (OutputRegister_n_65), .A (Product[1]), .B (\OutputRegister_register[1] ), .S (hfn_ipo_n72));
MUX2_X1 i_0_1_93 (.Z (OutputRegister_n_64), .A (Product[2]), .B (\OutputRegister_register[2] ), .S (hfn_ipo_n72));
MUX2_X1 i_0_1_92 (.Z (OutputRegister_n_63), .A (Product[3]), .B (\OutputRegister_register[3] ), .S (hfn_ipo_n72));
MUX2_X1 i_0_1_91 (.Z (OutputRegister_n_62), .A (Product[4]), .B (\OutputRegister_register[4] ), .S (hfn_ipo_n72));
MUX2_X1 i_0_1_90 (.Z (OutputRegister_n_61), .A (Product[5]), .B (\OutputRegister_register[5] ), .S (hfn_ipo_n72));
MUX2_X1 i_0_1_89 (.Z (OutputRegister_n_60), .A (Product[6]), .B (\OutputRegister_register[6] ), .S (hfn_ipo_n72));
MUX2_X1 i_0_1_88 (.Z (OutputRegister_n_59), .A (Product[7]), .B (\OutputRegister_register[7] ), .S (hfn_ipo_n72));
MUX2_X1 i_0_1_87 (.Z (OutputRegister_n_58), .A (Product[8]), .B (\OutputRegister_register[8] ), .S (hfn_ipo_n72));
MUX2_X1 i_0_1_86 (.Z (OutputRegister_n_57), .A (Product[9]), .B (\OutputRegister_register[9] ), .S (hfn_ipo_n72));
MUX2_X1 i_0_1_85 (.Z (OutputRegister_n_56), .A (Product[10]), .B (\OutputRegister_register[10] ), .S (hfn_ipo_n72));
MUX2_X1 i_0_1_84 (.Z (OutputRegister_n_55), .A (Product[11]), .B (\OutputRegister_register[11] ), .S (hfn_ipo_n72));
MUX2_X1 i_0_1_83 (.Z (OutputRegister_n_54), .A (Product[12]), .B (\OutputRegister_register[12] ), .S (enableA));
MUX2_X1 i_0_1_82 (.Z (OutputRegister_n_53), .A (Product[13]), .B (\OutputRegister_register[13] ), .S (enableA));
MUX2_X1 i_0_1_81 (.Z (OutputRegister_n_52), .A (Product[14]), .B (\OutputRegister_register[14] ), .S (enableA));
MUX2_X1 i_0_1_80 (.Z (OutputRegister_n_51), .A (Product[15]), .B (\OutputRegister_register[15] ), .S (enableA));
MUX2_X1 i_0_1_79 (.Z (OutputRegister_n_50), .A (Product[16]), .B (\OutputRegister_register[16] ), .S (enableA));
MUX2_X1 i_0_1_78 (.Z (OutputRegister_n_49), .A (Product[17]), .B (\OutputRegister_register[17] ), .S (enableA));
MUX2_X1 i_0_1_77 (.Z (OutputRegister_n_48), .A (Product[18]), .B (\OutputRegister_register[18] ), .S (enableA));
MUX2_X1 i_0_1_76 (.Z (OutputRegister_n_47), .A (Product[19]), .B (\OutputRegister_register[19] ), .S (enableA));
MUX2_X1 i_0_1_75 (.Z (OutputRegister_n_46), .A (Product[20]), .B (\OutputRegister_register[20] ), .S (enableA));
MUX2_X1 i_0_1_74 (.Z (OutputRegister_n_45), .A (Product[21]), .B (\OutputRegister_register[21] ), .S (enableA));
MUX2_X1 i_0_1_73 (.Z (OutputRegister_n_44), .A (Product[22]), .B (\OutputRegister_register[22] ), .S (hfn_ipo_n71));
MUX2_X1 i_0_1_72 (.Z (OutputRegister_n_43), .A (Product[23]), .B (\OutputRegister_register[23] ), .S (hfn_ipo_n71));
MUX2_X1 i_0_1_71 (.Z (OutputRegister_n_42), .A (Product[24]), .B (\OutputRegister_register[24] ), .S (hfn_ipo_n71));
MUX2_X1 i_0_1_70 (.Z (OutputRegister_n_41), .A (Product[25]), .B (\OutputRegister_register[25] ), .S (hfn_ipo_n71));
MUX2_X1 i_0_1_69 (.Z (OutputRegister_n_40), .A (Product[26]), .B (\OutputRegister_register[26] ), .S (hfn_ipo_n71));
MUX2_X1 i_0_1_68 (.Z (OutputRegister_n_39), .A (Product[27]), .B (\OutputRegister_register[27] ), .S (hfn_ipo_n71));
MUX2_X1 i_0_1_67 (.Z (OutputRegister_n_38), .A (Product[28]), .B (\OutputRegister_register[28] ), .S (hfn_ipo_n71));
MUX2_X1 i_0_1_66 (.Z (OutputRegister_n_37), .A (Product[29]), .B (\OutputRegister_register[29] ), .S (hfn_ipo_n71));
MUX2_X1 i_0_1_65 (.Z (OutputRegister_n_36), .A (Product[30]), .B (\OutputRegister_register[30] ), .S (hfn_ipo_n71));
MUX2_X1 i_0_1_64 (.Z (OutputRegister_n_35), .A (Product[31]), .B (\OutputRegister_register[31] ), .S (hfn_ipo_n71));
MUX2_X1 i_0_1_63 (.Z (OutputRegister_n_34), .A (Product[32]), .B (\OutputRegister_register[32] ), .S (hfn_ipo_n71));
MUX2_X1 i_0_1_62 (.Z (OutputRegister_n_33), .A (Product[33]), .B (\OutputRegister_register[33] ), .S (hfn_ipo_n71));
MUX2_X1 i_0_1_61 (.Z (OutputRegister_n_32), .A (Product[34]), .B (\OutputRegister_register[34] ), .S (hfn_ipo_n71));
MUX2_X1 i_0_1_60 (.Z (OutputRegister_n_31), .A (Product[35]), .B (\OutputRegister_register[35] ), .S (hfn_ipo_n71));
MUX2_X1 i_0_1_59 (.Z (OutputRegister_n_30), .A (Product[36]), .B (\OutputRegister_register[36] ), .S (hfn_ipo_n71));
MUX2_X1 i_0_1_58 (.Z (OutputRegister_n_29), .A (Product[37]), .B (\OutputRegister_register[37] ), .S (hfn_ipo_n71));
MUX2_X1 i_0_1_57 (.Z (OutputRegister_n_28), .A (Product[38]), .B (\OutputRegister_register[38] ), .S (hfn_ipo_n71));
MUX2_X1 i_0_1_56 (.Z (OutputRegister_n_27), .A (Product[39]), .B (\OutputRegister_register[39] ), .S (hfn_ipo_n71));
MUX2_X1 i_0_1_55 (.Z (OutputRegister_n_26), .A (Product[40]), .B (\OutputRegister_register[40] ), .S (hfn_ipo_n71));
MUX2_X1 i_0_1_54 (.Z (OutputRegister_n_25), .A (Product[41]), .B (\OutputRegister_register[41] ), .S (hfn_ipo_n71));
MUX2_X1 i_0_1_53 (.Z (OutputRegister_n_24), .A (Product[42]), .B (\OutputRegister_register[42] ), .S (hfn_ipo_n71));
MUX2_X1 i_0_1_52 (.Z (OutputRegister_n_23), .A (Product[43]), .B (\OutputRegister_register[43] ), .S (hfn_ipo_n71));
MUX2_X1 i_0_1_51 (.Z (OutputRegister_n_22), .A (Product[44]), .B (\OutputRegister_register[44] ), .S (hfn_ipo_n71));
MUX2_X1 i_0_1_50 (.Z (OutputRegister_n_21), .A (Product[45]), .B (\OutputRegister_register[45] ), .S (hfn_ipo_n71));
MUX2_X1 i_0_1_49 (.Z (OutputRegister_n_20), .A (Product[46]), .B (\OutputRegister_register[46] ), .S (hfn_ipo_n71));
MUX2_X1 i_0_1_48 (.Z (OutputRegister_n_19), .A (Product[47]), .B (\OutputRegister_register[47] ), .S (hfn_ipo_n71));
MUX2_X1 i_0_1_47 (.Z (OutputRegister_n_18), .A (Product[48]), .B (\OutputRegister_register[48] ), .S (hfn_ipo_n71));
MUX2_X1 i_0_1_46 (.Z (OutputRegister_n_17), .A (Product[49]), .B (\OutputRegister_register[49] ), .S (hfn_ipo_n71));
MUX2_X1 i_0_1_45 (.Z (OutputRegister_n_16), .A (Product[50]), .B (\OutputRegister_register[50] ), .S (hfn_ipo_n71));
MUX2_X1 i_0_1_44 (.Z (OutputRegister_n_15), .A (Product[51]), .B (\OutputRegister_register[51] ), .S (hfn_ipo_n71));
MUX2_X1 i_0_1_43 (.Z (OutputRegister_n_14), .A (Product[52]), .B (\OutputRegister_register[52] ), .S (hfn_ipo_n71));
MUX2_X1 i_0_1_42 (.Z (OutputRegister_n_13), .A (Product[53]), .B (\OutputRegister_register[53] ), .S (hfn_ipo_n71));
MUX2_X1 i_0_1_41 (.Z (OutputRegister_n_12), .A (Product[54]), .B (\OutputRegister_register[54] ), .S (hfn_ipo_n71));
MUX2_X1 i_0_1_40 (.Z (OutputRegister_n_11), .A (Product[55]), .B (\OutputRegister_register[55] ), .S (hfn_ipo_n71));
MUX2_X1 i_0_1_39 (.Z (OutputRegister_n_10), .A (Product[56]), .B (\OutputRegister_register[56] ), .S (hfn_ipo_n71));
MUX2_X1 i_0_1_38 (.Z (OutputRegister_n_9), .A (Product[57]), .B (\OutputRegister_register[57] ), .S (hfn_ipo_n71));
MUX2_X1 i_0_1_37 (.Z (OutputRegister_n_8), .A (Product[58]), .B (\OutputRegister_register[58] ), .S (hfn_ipo_n71));
MUX2_X1 i_0_1_36 (.Z (OutputRegister_n_7), .A (Product[59]), .B (\OutputRegister_register[59] ), .S (hfn_ipo_n71));
MUX2_X1 i_0_1_35 (.Z (OutputRegister_n_6), .A (Product[60]), .B (\OutputRegister_register[60] ), .S (hfn_ipo_n71));
MUX2_X1 i_0_1_34 (.Z (OutputRegister_n_5), .A (Product[61]), .B (\OutputRegister_register[61] ), .S (hfn_ipo_n71));
MUX2_X1 i_0_1_33 (.Z (OutputRegister_n_4), .A (Product[62]), .B (\OutputRegister_register[62] ), .S (hfn_ipo_n71));
MUX2_X1 i_0_1_32 (.Z (OutputRegister_n_2), .A (Product[63]), .B (\OutputRegister_register[63] ), .S (hfn_ipo_n71));
MUX2_X1 i_0_1_31 (.Z (InputRegisterA_n_34), .A (slo__n236), .B (\InputRegisterA_register[0] ), .S (hfn_ipo_n72));
MUX2_X1 i_0_1_30 (.Z (InputRegisterA_n_33), .A (slo__n198), .B (\InputRegisterA_register[1] ), .S (hfn_ipo_n72));
MUX2_X1 i_0_1_29 (.Z (InputRegisterA_n_32), .A (\registerOutA[2] ), .B (\InputRegisterA_register[2] ), .S (hfn_ipo_n72));
MUX2_X1 i_0_1_28 (.Z (InputRegisterA_n_31), .A (\registerOutA[3] ), .B (\InputRegisterA_register[3] ), .S (hfn_ipo_n72));
MUX2_X1 i_0_1_27 (.Z (InputRegisterA_n_30), .A (\registerOutA[4] ), .B (\InputRegisterA_register[4] ), .S (hfn_ipo_n72));
MUX2_X1 i_0_1_26 (.Z (InputRegisterA_n_29), .A (\registerOutA[5] ), .B (\InputRegisterA_register[5] ), .S (hfn_ipo_n72));
MUX2_X1 i_0_1_25 (.Z (InputRegisterA_n_28), .A (\registerOutA[6] ), .B (\InputRegisterA_register[6] ), .S (hfn_ipo_n72));
MUX2_X1 i_0_1_24 (.Z (InputRegisterA_n_27), .A (\registerOutA[7] ), .B (\InputRegisterA_register[7] ), .S (hfn_ipo_n72));
MUX2_X1 i_0_1_23 (.Z (InputRegisterA_n_26), .A (\registerOutA[8] ), .B (\InputRegisterA_register[8] ), .S (hfn_ipo_n72));
MUX2_X1 i_0_1_22 (.Z (InputRegisterA_n_25), .A (\registerOutA[9] ), .B (\InputRegisterA_register[9] ), .S (hfn_ipo_n72));
MUX2_X1 i_0_1_21 (.Z (InputRegisterA_n_24), .A (\registerOutA[10] ), .B (\InputRegisterA_register[10] ), .S (hfn_ipo_n72));
MUX2_X1 i_0_1_20 (.Z (InputRegisterA_n_23), .A (\registerOutA[11] ), .B (\InputRegisterA_register[11] ), .S (hfn_ipo_n72));
MUX2_X1 i_0_1_19 (.Z (InputRegisterA_n_22), .A (\registerOutA[12] ), .B (\InputRegisterA_register[12] ), .S (hfn_ipo_n72));
MUX2_X1 i_0_1_18 (.Z (InputRegisterA_n_21), .A (\registerOutA[13] ), .B (\InputRegisterA_register[13] ), .S (hfn_ipo_n72));
MUX2_X1 i_0_1_17 (.Z (InputRegisterA_n_20), .A (\registerOutA[14] ), .B (\InputRegisterA_register[14] ), .S (enableA));
MUX2_X1 i_0_1_16 (.Z (InputRegisterA_n_19), .A (\registerOutA[15] ), .B (\InputRegisterA_register[15] ), .S (hfn_ipo_n72));
MUX2_X1 i_0_1_15 (.Z (InputRegisterA_n_18), .A (\registerOutA[16] ), .B (\InputRegisterA_register[16] ), .S (enableA));
MUX2_X1 i_0_1_14 (.Z (InputRegisterA_n_17), .A (\registerOutA[17] ), .B (\InputRegisterA_register[17] ), .S (enableA));
MUX2_X1 i_0_1_13 (.Z (InputRegisterA_n_16), .A (\registerOutA[18] ), .B (\InputRegisterA_register[18] ), .S (enableA));
MUX2_X1 i_0_1_12 (.Z (InputRegisterA_n_15), .A (\registerOutA[19] ), .B (\InputRegisterA_register[19] ), .S (enableA));
MUX2_X1 i_0_1_11 (.Z (InputRegisterA_n_14), .A (\registerOutA[20] ), .B (\InputRegisterA_register[20] ), .S (enableA));
MUX2_X1 i_0_1_10 (.Z (InputRegisterA_n_13), .A (\registerOutA[21] ), .B (\InputRegisterA_register[21] ), .S (enableA));
MUX2_X1 i_0_1_9 (.Z (InputRegisterA_n_12), .A (\registerOutA[22] ), .B (\InputRegisterA_register[22] ), .S (enableA));
MUX2_X1 i_0_1_8 (.Z (InputRegisterA_n_11), .A (\registerOutA[23] ), .B (\InputRegisterA_register[23] ), .S (enableA));
MUX2_X1 i_0_1_7 (.Z (InputRegisterA_n_10), .A (\registerOutA[24] ), .B (\InputRegisterA_register[24] ), .S (enableA));
MUX2_X1 i_0_1_6 (.Z (InputRegisterA_n_9), .A (\registerOutA[25] ), .B (\InputRegisterA_register[25] ), .S (hfn_ipo_n71));
MUX2_X1 i_0_1_5 (.Z (InputRegisterA_n_8), .A (\registerOutA[26] ), .B (\InputRegisterA_register[26] ), .S (hfn_ipo_n71));
MUX2_X1 i_0_1_4 (.Z (InputRegisterA_n_7), .A (\registerOutA[27] ), .B (\InputRegisterA_register[27] ), .S (hfn_ipo_n71));
MUX2_X1 i_0_1_3 (.Z (InputRegisterA_n_6), .A (\registerOutA[28] ), .B (\InputRegisterA_register[28] ), .S (hfn_ipo_n72));
MUX2_X1 i_0_1_2 (.Z (InputRegisterA_n_5), .A (\registerOutA[29] ), .B (\InputRegisterA_register[29] ), .S (hfn_ipo_n72));
MUX2_X1 i_0_1_1 (.Z (InputRegisterA_n_4), .A (\registerOutA[30] ), .B (\InputRegisterA_register[30] ), .S (hfn_ipo_n72));
MUX2_X1 i_0_1_0 (.Z (InputRegisterA_n_2), .A (\registerOutA[31] ), .B (\InputRegisterA_register[31] ), .S (hfn_ipo_n72));
MUX2_X1 i_0_0_31 (.Z (InputRegisterB_n_34), .A (opt_ipo_n299), .B (\InputRegisterB_register[0] ), .S (enableB));
MUX2_X1 i_0_0_30 (.Z (InputRegisterB_n_33), .A (drc_ipo_n76), .B (\InputRegisterB_register[1] ), .S (enableB));
MUX2_X1 i_0_0_29 (.Z (InputRegisterB_n_32), .A (\registerOutB[2] ), .B (\InputRegisterB_register[2] ), .S (enableB));
MUX2_X1 i_0_0_28 (.Z (InputRegisterB_n_31), .A (drc_ipo_n78), .B (\InputRegisterB_register[3] ), .S (enableB));
MUX2_X1 i_0_0_27 (.Z (InputRegisterB_n_30), .A (drc_ipo_n79), .B (\InputRegisterB_register[4] ), .S (enableB));
MUX2_X1 i_0_0_26 (.Z (InputRegisterB_n_29), .A (drc_ipo_n80), .B (\InputRegisterB_register[5] ), .S (enableB));
MUX2_X1 i_0_0_25 (.Z (InputRegisterB_n_28), .A (\registerOutB[6] ), .B (\InputRegisterB_register[6] ), .S (enableB));
MUX2_X1 i_0_0_24 (.Z (InputRegisterB_n_27), .A (drc_ipo_n82), .B (\InputRegisterB_register[7] ), .S (enableB));
MUX2_X1 i_0_0_23 (.Z (InputRegisterB_n_26), .A (drc_ipo_n347), .B (\InputRegisterB_register[8] ), .S (enableB));
MUX2_X1 i_0_0_22 (.Z (InputRegisterB_n_25), .A (drc_ipo_n348), .B (\InputRegisterB_register[9] ), .S (enableB));
MUX2_X1 i_0_0_21 (.Z (InputRegisterB_n_24), .A (drc_ipo_n85), .B (\InputRegisterB_register[10] ), .S (enableB));
MUX2_X1 i_0_0_20 (.Z (InputRegisterB_n_23), .A (drc_ipo_n86), .B (\InputRegisterB_register[11] ), .S (enableB));
MUX2_X1 i_0_0_19 (.Z (InputRegisterB_n_22), .A (drc_ipo_n87), .B (\InputRegisterB_register[12] ), .S (enableB));
MUX2_X1 i_0_0_18 (.Z (InputRegisterB_n_21), .A (drc_ipo_n88), .B (\InputRegisterB_register[13] ), .S (enableB));
MUX2_X1 i_0_0_17 (.Z (InputRegisterB_n_20), .A (drc_ipo_n89), .B (\InputRegisterB_register[14] ), .S (enableB));
MUX2_X1 i_0_0_16 (.Z (InputRegisterB_n_19), .A (drc_ipo_n90), .B (\InputRegisterB_register[15] ), .S (enableB));
MUX2_X1 i_0_0_15 (.Z (InputRegisterB_n_18), .A (drc_ipo_n350), .B (\InputRegisterB_register[16] ), .S (enableB));
MUX2_X1 i_0_0_14 (.Z (InputRegisterB_n_17), .A (drc_ipo_n351), .B (\InputRegisterB_register[17] ), .S (enableB));
MUX2_X1 i_0_0_13 (.Z (InputRegisterB_n_16), .A (drc_ipo_n93), .B (\InputRegisterB_register[18] ), .S (enableB));
MUX2_X1 i_0_0_12 (.Z (InputRegisterB_n_15), .A (drc_ipo_n94), .B (\InputRegisterB_register[19] ), .S (enableB));
MUX2_X1 i_0_0_11 (.Z (InputRegisterB_n_14), .A (drc_ipo_n95), .B (\InputRegisterB_register[20] ), .S (enableB));
MUX2_X1 i_0_0_10 (.Z (InputRegisterB_n_13), .A (drc_ipo_n96), .B (\InputRegisterB_register[21] ), .S (enableB));
MUX2_X1 i_0_0_9 (.Z (InputRegisterB_n_12), .A (drc_ipo_n97), .B (\InputRegisterB_register[22] ), .S (enableB));
MUX2_X1 i_0_0_8 (.Z (InputRegisterB_n_11), .A (drc_ipo_n352), .B (\InputRegisterB_register[23] ), .S (enableB));
MUX2_X1 i_0_0_7 (.Z (InputRegisterB_n_10), .A (drc_ipo_n99), .B (\InputRegisterB_register[24] ), .S (enableB));
MUX2_X1 i_0_0_6 (.Z (InputRegisterB_n_9), .A (drc_ipo_n100), .B (\InputRegisterB_register[25] ), .S (enableB));
MUX2_X1 i_0_0_5 (.Z (InputRegisterB_n_8), .A (drc_ipo_n353), .B (\InputRegisterB_register[26] ), .S (enableB));
MUX2_X1 i_0_0_4 (.Z (InputRegisterB_n_7), .A (drc_ipo_n355), .B (\InputRegisterB_register[27] ), .S (enableB));
MUX2_X1 i_0_0_3 (.Z (InputRegisterB_n_6), .A (drc_ipo_n103), .B (\InputRegisterB_register[28] ), .S (enableB));
MUX2_X1 i_0_0_2 (.Z (InputRegisterB_n_5), .A (drc_ipo_n104), .B (\InputRegisterB_register[29] ), .S (enableB));
MUX2_X1 i_0_0_1 (.Z (InputRegisterB_n_4), .A (\registerOutB[30] ), .B (\InputRegisterB_register[30] ), .S (enableB));
MUX2_X1 i_0_0_0 (.Z (InputRegisterB_n_2), .A (drc_ipo_n105), .B (\InputRegisterB_register[31] ), .S (enableB));
INV_X16 CTS_L6_c609 (.ZN (CTS_n617), .A (CTS_n630));
INV_X1 OutputRegister_i_0_0 (.ZN (OutputRegister_n_1), .A (resetOut));
INV_X2 InputRegisterB_i_0_0 (.ZN (InputRegisterB_n_1), .A (resetB));
INV_X2 InputRegisterA_i_0_0 (.ZN (InputRegisterA_n_1), .A (resetA));
DFF_X1 \OutputRegister_dataOut_reg[0]  (.Q (Product[0]), .CK (CTS_n618), .D (OutputRegister_n_66));
DFF_X1 \OutputRegister_dataOut_reg[1]  (.Q (Product[1]), .CK (CTS_n618), .D (OutputRegister_n_65));
DFF_X1 \OutputRegister_dataOut_reg[2]  (.Q (Product[2]), .CK (CTS_n618), .D (OutputRegister_n_64));
DFF_X1 \OutputRegister_dataOut_reg[3]  (.Q (Product[3]), .CK (CTS_n618), .D (OutputRegister_n_63));
DFF_X1 \OutputRegister_dataOut_reg[4]  (.Q (Product[4]), .CK (CTS_n618), .D (OutputRegister_n_62));
DFF_X1 \OutputRegister_dataOut_reg[5]  (.Q (Product[5]), .CK (CTS_n618), .D (OutputRegister_n_61));
DFF_X1 \OutputRegister_dataOut_reg[6]  (.Q (Product[6]), .CK (CTS_n618), .D (OutputRegister_n_60));
DFF_X1 \OutputRegister_dataOut_reg[7]  (.Q (Product[7]), .CK (CTS_n618), .D (OutputRegister_n_59));
DFF_X1 \OutputRegister_dataOut_reg[8]  (.Q (Product[8]), .CK (CTS_n618), .D (OutputRegister_n_58));
DFF_X1 \OutputRegister_dataOut_reg[9]  (.Q (Product[9]), .CK (CTS_n618), .D (OutputRegister_n_57));
DFF_X1 \OutputRegister_dataOut_reg[10]  (.Q (Product[10]), .CK (CTS_n617), .D (OutputRegister_n_56));
DFF_X1 \OutputRegister_dataOut_reg[11]  (.Q (Product[11]), .CK (CTS_n617), .D (OutputRegister_n_55));
DFF_X1 \OutputRegister_dataOut_reg[12]  (.Q (Product[12]), .CK (CTS_n617), .D (OutputRegister_n_54));
DFF_X1 \OutputRegister_dataOut_reg[13]  (.Q (Product[13]), .CK (CTS_n617), .D (OutputRegister_n_53));
DFF_X1 \OutputRegister_dataOut_reg[14]  (.Q (Product[14]), .CK (CTS_n617), .D (OutputRegister_n_52));
DFF_X1 \OutputRegister_dataOut_reg[15]  (.Q (Product[15]), .CK (CTS_n617), .D (OutputRegister_n_51));
DFF_X1 \OutputRegister_dataOut_reg[16]  (.Q (Product[16]), .CK (CTS_n617), .D (OutputRegister_n_50));
DFF_X1 \OutputRegister_dataOut_reg[17]  (.Q (Product[17]), .CK (CTS_n617), .D (OutputRegister_n_49));
DFF_X1 \OutputRegister_dataOut_reg[18]  (.Q (Product[18]), .CK (CTS_n617), .D (OutputRegister_n_48));
DFF_X1 \OutputRegister_dataOut_reg[19]  (.Q (Product[19]), .CK (CTS_n617), .D (OutputRegister_n_47));
DFF_X1 \OutputRegister_dataOut_reg[20]  (.Q (Product[20]), .CK (CTS_n617), .D (OutputRegister_n_46));
DFF_X1 \OutputRegister_dataOut_reg[21]  (.Q (Product[21]), .CK (CTS_n617), .D (OutputRegister_n_45));
DFF_X1 \OutputRegister_dataOut_reg[22]  (.Q (Product[22]), .CK (CTS_n619), .D (OutputRegister_n_44));
DFF_X1 \OutputRegister_dataOut_reg[23]  (.Q (Product[23]), .CK (CTS_n619), .D (OutputRegister_n_43));
DFF_X1 \OutputRegister_dataOut_reg[24]  (.Q (Product[24]), .CK (CTS_n619), .D (OutputRegister_n_42));
DFF_X1 \OutputRegister_dataOut_reg[25]  (.Q (Product[25]), .CK (CTS_n619), .D (OutputRegister_n_41));
DFF_X1 \OutputRegister_dataOut_reg[26]  (.Q (Product[26]), .CK (CTS_n619), .D (OutputRegister_n_40));
DFF_X1 \OutputRegister_dataOut_reg[27]  (.Q (Product[27]), .CK (CTS_n619), .D (OutputRegister_n_39));
DFF_X1 \OutputRegister_dataOut_reg[28]  (.Q (Product[28]), .CK (CTS_n619), .D (OutputRegister_n_38));
DFF_X1 \OutputRegister_dataOut_reg[29]  (.Q (Product[29]), .CK (CTS_n619), .D (OutputRegister_n_37));
DFF_X1 \OutputRegister_dataOut_reg[30]  (.Q (Product[30]), .CK (CTS_n619), .D (OutputRegister_n_36));
DFF_X1 \OutputRegister_dataOut_reg[31]  (.Q (Product[31]), .CK (CTS_n619), .D (OutputRegister_n_35));
DFF_X1 \OutputRegister_dataOut_reg[32]  (.Q (Product[32]), .CK (CTS_n619), .D (OutputRegister_n_34));
DFF_X1 \OutputRegister_dataOut_reg[33]  (.Q (Product[33]), .CK (CTS_n619), .D (OutputRegister_n_33));
DFF_X1 \OutputRegister_dataOut_reg[34]  (.Q (Product[34]), .CK (CTS_n619), .D (OutputRegister_n_32));
DFF_X1 \OutputRegister_dataOut_reg[35]  (.Q (Product[35]), .CK (CTS_n619), .D (OutputRegister_n_31));
DFF_X1 \OutputRegister_dataOut_reg[36]  (.Q (Product[36]), .CK (CTS_n619), .D (OutputRegister_n_30));
DFF_X1 \OutputRegister_dataOut_reg[37]  (.Q (Product[37]), .CK (CTS_n619), .D (OutputRegister_n_29));
DFF_X1 \OutputRegister_dataOut_reg[38]  (.Q (Product[38]), .CK (CTS_n619), .D (OutputRegister_n_28));
DFF_X1 \OutputRegister_dataOut_reg[39]  (.Q (Product[39]), .CK (CTS_n619), .D (OutputRegister_n_27));
DFF_X1 \OutputRegister_dataOut_reg[40]  (.Q (Product[40]), .CK (CTS_n619), .D (OutputRegister_n_26));
DFF_X1 \OutputRegister_dataOut_reg[41]  (.Q (Product[41]), .CK (CTS_n619), .D (OutputRegister_n_25));
DFF_X1 \OutputRegister_dataOut_reg[42]  (.Q (Product[42]), .CK (CTS_n619), .D (OutputRegister_n_24));
DFF_X1 \OutputRegister_dataOut_reg[43]  (.Q (Product[43]), .CK (CTS_n619), .D (OutputRegister_n_23));
DFF_X1 \OutputRegister_dataOut_reg[44]  (.Q (Product[44]), .CK (CTS_n619), .D (OutputRegister_n_22));
DFF_X1 \OutputRegister_dataOut_reg[45]  (.Q (Product[45]), .CK (CTS_n619), .D (OutputRegister_n_21));
DFF_X1 \OutputRegister_dataOut_reg[46]  (.Q (Product[46]), .CK (CTS_n619), .D (OutputRegister_n_20));
DFF_X1 \OutputRegister_dataOut_reg[47]  (.Q (Product[47]), .CK (CTS_n619), .D (OutputRegister_n_19));
DFF_X1 \OutputRegister_dataOut_reg[48]  (.Q (Product[48]), .CK (CTS_n619), .D (OutputRegister_n_18));
DFF_X1 \OutputRegister_dataOut_reg[49]  (.Q (Product[49]), .CK (CTS_n619), .D (OutputRegister_n_17));
DFF_X1 \OutputRegister_dataOut_reg[50]  (.Q (Product[50]), .CK (CTS_n619), .D (OutputRegister_n_16));
DFF_X1 \OutputRegister_dataOut_reg[51]  (.Q (Product[51]), .CK (CTS_n619), .D (OutputRegister_n_15));
DFF_X1 \OutputRegister_dataOut_reg[52]  (.Q (Product[52]), .CK (CTS_n619), .D (OutputRegister_n_14));
DFF_X1 \OutputRegister_dataOut_reg[53]  (.Q (Product[53]), .CK (CTS_n619), .D (OutputRegister_n_13));
DFF_X1 \OutputRegister_dataOut_reg[54]  (.Q (Product[54]), .CK (CTS_n619), .D (OutputRegister_n_12));
DFF_X1 \OutputRegister_dataOut_reg[55]  (.Q (Product[55]), .CK (CTS_n618), .D (OutputRegister_n_11));
DFF_X1 \OutputRegister_dataOut_reg[56]  (.Q (Product[56]), .CK (CTS_n619), .D (OutputRegister_n_10));
DFF_X1 \OutputRegister_dataOut_reg[57]  (.Q (Product[57]), .CK (CTS_n619), .D (OutputRegister_n_9));
DFF_X1 \OutputRegister_dataOut_reg[58]  (.Q (Product[58]), .CK (CTS_n619), .D (OutputRegister_n_8));
DFF_X1 \OutputRegister_dataOut_reg[59]  (.Q (Product[59]), .CK (CTS_n619), .D (OutputRegister_n_7));
DFF_X1 \OutputRegister_dataOut_reg[60]  (.Q (Product[60]), .CK (CTS_n619), .D (OutputRegister_n_6));
DFF_X1 \OutputRegister_dataOut_reg[61]  (.Q (Product[61]), .CK (CTS_n619), .D (OutputRegister_n_5));
DFF_X1 \OutputRegister_dataOut_reg[62]  (.Q (Product[62]), .CK (CTS_n619), .D (OutputRegister_n_4));
DFF_X1 \OutputRegister_dataOut_reg[63]  (.Q (Product[63]), .CK (CTS_n619), .D (OutputRegister_n_2));
DFFR_X1 \OutputRegister_register_reg[0]  (.Q (\OutputRegister_register[0] ), .CK (CTS_n564)
    , .D (\registerInProduct[0] ), .RN (hfn_ipo_n74));
DFFR_X1 \OutputRegister_register_reg[1]  (.Q (\OutputRegister_register[1] ), .CK (CTS_n564)
    , .D (\registerInProduct[1] ), .RN (hfn_ipo_n74));
DFFR_X1 \OutputRegister_register_reg[2]  (.Q (\OutputRegister_register[2] ), .CK (CTS_n564)
    , .D (\registerInProduct[2] ), .RN (hfn_ipo_n74));
DFFR_X1 \OutputRegister_register_reg[3]  (.Q (\OutputRegister_register[3] ), .CK (CTS_n564)
    , .D (\registerInProduct[3] ), .RN (hfn_ipo_n74));
DFFR_X1 \OutputRegister_register_reg[4]  (.Q (\OutputRegister_register[4] ), .CK (CTS_n564)
    , .D (\registerInProduct[4] ), .RN (hfn_ipo_n74));
DFFR_X1 \OutputRegister_register_reg[5]  (.Q (\OutputRegister_register[5] ), .CK (CTS_n564)
    , .D (\registerInProduct[5] ), .RN (hfn_ipo_n74));
DFFR_X1 \OutputRegister_register_reg[6]  (.Q (\OutputRegister_register[6] ), .CK (CTS_n564)
    , .D (\registerInProduct[6] ), .RN (hfn_ipo_n74));
DFFR_X1 \OutputRegister_register_reg[7]  (.Q (\OutputRegister_register[7] ), .CK (CTS_n564)
    , .D (\registerInProduct[7] ), .RN (hfn_ipo_n74));
DFFR_X1 \OutputRegister_register_reg[8]  (.Q (\OutputRegister_register[8] ), .CK (CTS_n564)
    , .D (\registerInProduct[8] ), .RN (hfn_ipo_n74));
DFFR_X1 \OutputRegister_register_reg[9]  (.Q (\OutputRegister_register[9] ), .CK (CTS_n564)
    , .D (\registerInProduct[9] ), .RN (hfn_ipo_n74));
DFFR_X1 \OutputRegister_register_reg[10]  (.Q (\OutputRegister_register[10] ), .CK (CTS_n564)
    , .D (\registerInProduct[10] ), .RN (CLOCK_spc__n1018));
DFFR_X1 \OutputRegister_register_reg[11]  (.Q (\OutputRegister_register[11] ), .CK (CTS_n564)
    , .D (\registerInProduct[11] ), .RN (CLOCK_spc__n1018));
DFFR_X1 \OutputRegister_register_reg[12]  (.Q (\OutputRegister_register[12] ), .CK (CTS_n564)
    , .D (\registerInProduct[12] ), .RN (CLOCK_spc__n1018));
DFFR_X1 \OutputRegister_register_reg[13]  (.Q (\OutputRegister_register[13] ), .CK (CTS_n564)
    , .D (\registerInProduct[13] ), .RN (CLOCK_spc__n1018));
DFFR_X1 \OutputRegister_register_reg[14]  (.Q (\OutputRegister_register[14] ), .CK (CTS_n564)
    , .D (\registerInProduct[14] ), .RN (CLOCK_spc__n1018));
DFFR_X1 \OutputRegister_register_reg[15]  (.Q (\OutputRegister_register[15] ), .CK (CTS_n564)
    , .D (\registerInProduct[15] ), .RN (CLOCK_spc__n1018));
DFFR_X1 \OutputRegister_register_reg[16]  (.Q (\OutputRegister_register[16] ), .CK (CTS_n564)
    , .D (\registerInProduct[16] ), .RN (CLOCK_spc__n1018));
DFFR_X1 \OutputRegister_register_reg[17]  (.Q (\OutputRegister_register[17] ), .CK (CTS_n564)
    , .D (\registerInProduct[17] ), .RN (CLOCK_spc__n1018));
DFFR_X1 \OutputRegister_register_reg[18]  (.Q (\OutputRegister_register[18] ), .CK (CTS_n564)
    , .D (\registerInProduct[18] ), .RN (CLOCK_spc__n1018));
DFFR_X1 \OutputRegister_register_reg[19]  (.Q (\OutputRegister_register[19] ), .CK (CTS_n564)
    , .D (\registerInProduct[19] ), .RN (CLOCK_spc__n1018));
DFFR_X1 \OutputRegister_register_reg[20]  (.Q (\OutputRegister_register[20] ), .CK (CTS_n564)
    , .D (\registerInProduct[20] ), .RN (CLOCK_spc__n1018));
DFFR_X1 \OutputRegister_register_reg[21]  (.Q (\OutputRegister_register[21] ), .CK (CTS_n564)
    , .D (\registerInProduct[21] ), .RN (CLOCK_spc__n1018));
DFFR_X1 \OutputRegister_register_reg[22]  (.Q (\OutputRegister_register[22] ), .CK (CTS_n565)
    , .D (\registerInProduct[22] ), .RN (CLOCK_spc__n1018));
DFFR_X1 \OutputRegister_register_reg[23]  (.Q (\OutputRegister_register[23] ), .CK (CTS_n565)
    , .D (\registerInProduct[23] ), .RN (CLOCK_spc__n1018));
DFFR_X1 \OutputRegister_register_reg[24]  (.Q (\OutputRegister_register[24] ), .CK (CTS_n565)
    , .D (\registerInProduct[24] ), .RN (CLOCK_spc__n1018));
DFFR_X1 \OutputRegister_register_reg[25]  (.Q (\OutputRegister_register[25] ), .CK (CTS_n565)
    , .D (\registerInProduct[25] ), .RN (CLOCK_spc__n1018));
DFFR_X1 \OutputRegister_register_reg[26]  (.Q (\OutputRegister_register[26] ), .CK (CTS_n565)
    , .D (\registerInProduct[26] ), .RN (CLOCK_spc__n1018));
DFFR_X1 \OutputRegister_register_reg[27]  (.Q (\OutputRegister_register[27] ), .CK (CTS_n565)
    , .D (\registerInProduct[27] ), .RN (CLOCK_spc__n1018));
DFFR_X1 \OutputRegister_register_reg[28]  (.Q (\OutputRegister_register[28] ), .CK (CTS_n565)
    , .D (\registerInProduct[28] ), .RN (CLOCK_spc__n1018));
DFFR_X1 \OutputRegister_register_reg[29]  (.Q (\OutputRegister_register[29] ), .CK (CTS_n565)
    , .D (\registerInProduct[29] ), .RN (CLOCK_spc__n1018));
DFFR_X1 \OutputRegister_register_reg[30]  (.Q (\OutputRegister_register[30] ), .CK (CTS_n565)
    , .D (\registerInProduct[30] ), .RN (CLOCK_spc__n1018));
DFFR_X1 \OutputRegister_register_reg[31]  (.Q (\OutputRegister_register[31] ), .CK (CTS_n565)
    , .D (\registerInProduct[31] ), .RN (OutputRegister_n_1));
DFFR_X1 \OutputRegister_register_reg[32]  (.Q (\OutputRegister_register[32] ), .CK (CTS_n565)
    , .D (\registerInProduct[32] ), .RN (CLOCK_spc__n1018));
DFFR_X1 \OutputRegister_register_reg[33]  (.Q (\OutputRegister_register[33] ), .CK (CTS_n565)
    , .D (\registerInProduct[33] ), .RN (CLOCK_spc__n1018));
DFFR_X1 \OutputRegister_register_reg[34]  (.Q (\OutputRegister_register[34] ), .CK (CTS_n565)
    , .D (\registerInProduct[34] ), .RN (hfn_ipo_n74));
DFFR_X1 \OutputRegister_register_reg[35]  (.Q (\OutputRegister_register[35] ), .CK (CTS_n565)
    , .D (\registerInProduct[35] ), .RN (hfn_ipo_n74));
DFFR_X1 \OutputRegister_register_reg[36]  (.Q (\OutputRegister_register[36] ), .CK (CTS_n565)
    , .D (\registerInProduct[36] ), .RN (hfn_ipo_n74));
DFFR_X1 \OutputRegister_register_reg[37]  (.Q (\OutputRegister_register[37] ), .CK (CTS_n565)
    , .D (\registerInProduct[37] ), .RN (hfn_ipo_n74));
DFFR_X1 \OutputRegister_register_reg[38]  (.Q (\OutputRegister_register[38] ), .CK (CTS_n565)
    , .D (\registerInProduct[38] ), .RN (hfn_ipo_n74));
DFFR_X1 \OutputRegister_register_reg[39]  (.Q (\OutputRegister_register[39] ), .CK (CTS_n565)
    , .D (\registerInProduct[39] ), .RN (hfn_ipo_n74));
DFFR_X1 \OutputRegister_register_reg[40]  (.Q (\OutputRegister_register[40] ), .CK (CTS_n565)
    , .D (\registerInProduct[40] ), .RN (hfn_ipo_n74));
DFFR_X1 \OutputRegister_register_reg[41]  (.Q (\OutputRegister_register[41] ), .CK (CTS_n565)
    , .D (\registerInProduct[41] ), .RN (hfn_ipo_n74));
DFFR_X1 \OutputRegister_register_reg[42]  (.Q (\OutputRegister_register[42] ), .CK (CTS_n565)
    , .D (\registerInProduct[42] ), .RN (hfn_ipo_n74));
DFFR_X1 \OutputRegister_register_reg[43]  (.Q (\OutputRegister_register[43] ), .CK (CTS_n565)
    , .D (\registerInProduct[43] ), .RN (hfn_ipo_n74));
DFFR_X1 \OutputRegister_register_reg[44]  (.Q (\OutputRegister_register[44] ), .CK (CTS_n565)
    , .D (\registerInProduct[44] ), .RN (hfn_ipo_n74));
DFFR_X1 \OutputRegister_register_reg[45]  (.Q (\OutputRegister_register[45] ), .CK (CTS_n565)
    , .D (\registerInProduct[45] ), .RN (hfn_ipo_n74));
DFFR_X1 \OutputRegister_register_reg[46]  (.Q (\OutputRegister_register[46] ), .CK (CTS_n565)
    , .D (\registerInProduct[46] ), .RN (hfn_ipo_n74));
DFFR_X1 \OutputRegister_register_reg[47]  (.Q (\OutputRegister_register[47] ), .CK (CTS_n565)
    , .D (\registerInProduct[47] ), .RN (hfn_ipo_n74));
DFFR_X1 \OutputRegister_register_reg[48]  (.Q (\OutputRegister_register[48] ), .CK (CTS_n565)
    , .D (\registerInProduct[48] ), .RN (hfn_ipo_n74));
DFFR_X1 \OutputRegister_register_reg[49]  (.Q (\OutputRegister_register[49] ), .CK (CTS_n565)
    , .D (\registerInProduct[49] ), .RN (hfn_ipo_n74));
DFFR_X1 \OutputRegister_register_reg[50]  (.Q (\OutputRegister_register[50] ), .CK (CTS_n565)
    , .D (\registerInProduct[50] ), .RN (hfn_ipo_n74));
DFFR_X1 \OutputRegister_register_reg[51]  (.Q (\OutputRegister_register[51] ), .CK (CTS_n565)
    , .D (\registerInProduct[51] ), .RN (hfn_ipo_n74));
DFFR_X1 \OutputRegister_register_reg[52]  (.Q (\OutputRegister_register[52] ), .CK (CTS_n565)
    , .D (\registerInProduct[52] ), .RN (hfn_ipo_n74));
DFFR_X1 \OutputRegister_register_reg[53]  (.Q (\OutputRegister_register[53] ), .CK (CTS_n565)
    , .D (\registerInProduct[53] ), .RN (hfn_ipo_n74));
DFFR_X1 \OutputRegister_register_reg[54]  (.Q (\OutputRegister_register[54] ), .CK (CTS_n565)
    , .D (\registerInProduct[54] ), .RN (hfn_ipo_n74));
DFFR_X1 \OutputRegister_register_reg[55]  (.Q (\OutputRegister_register[55] ), .CK (CTS_n565)
    , .D (\registerInProduct[55] ), .RN (hfn_ipo_n74));
DFFR_X1 \OutputRegister_register_reg[56]  (.Q (\OutputRegister_register[56] ), .CK (CTS_n565)
    , .D (\registerInProduct[56] ), .RN (hfn_ipo_n74));
DFFR_X1 \OutputRegister_register_reg[57]  (.Q (\OutputRegister_register[57] ), .CK (CTS_n565)
    , .D (\registerInProduct[57] ), .RN (hfn_ipo_n74));
DFFR_X1 \OutputRegister_register_reg[58]  (.Q (\OutputRegister_register[58] ), .CK (CTS_n565)
    , .D (\registerInProduct[58] ), .RN (hfn_ipo_n74));
DFFR_X1 \OutputRegister_register_reg[59]  (.Q (\OutputRegister_register[59] ), .CK (CTS_n565)
    , .D (\registerInProduct[59] ), .RN (hfn_ipo_n74));
DFFR_X1 \OutputRegister_register_reg[60]  (.Q (\OutputRegister_register[60] ), .CK (CTS_n565)
    , .D (\registerInProduct[60] ), .RN (hfn_ipo_n74));
DFFR_X1 \OutputRegister_register_reg[61]  (.Q (\OutputRegister_register[61] ), .CK (CTS_n565)
    , .D (\registerInProduct[61] ), .RN (hfn_ipo_n74));
DFFR_X1 \OutputRegister_register_reg[62]  (.Q (\OutputRegister_register[62] ), .CK (CTS_n565)
    , .D (\registerInProduct[62] ), .RN (hfn_ipo_n74));
DFFR_X1 \OutputRegister_register_reg[63]  (.Q (\OutputRegister_register[63] ), .CK (CTS_n565)
    , .D (\registerInProduct[63] ), .RN (hfn_ipo_n74));
DFF_X1 \InputRegisterB_dataOut_reg[0]  (.Q (slo___n231), .CK (CTS_n617), .D (InputRegisterB_n_34));
DFF_X1 \InputRegisterB_dataOut_reg[1]  (.Q (\registerOutB[1] ), .CK (CTS_n617), .D (InputRegisterB_n_33));
DFF_X1 \InputRegisterB_dataOut_reg[2]  (.Q (\registerOutB[2] ), .CK (CTS_n617), .D (InputRegisterB_n_32));
DFF_X1 \InputRegisterB_dataOut_reg[3]  (.Q (\registerOutB[3] ), .CK (CTS_n618), .D (InputRegisterB_n_31));
DFF_X1 \InputRegisterB_dataOut_reg[4]  (.Q (\registerOutB[4] ), .CK (CTS_n617), .D (InputRegisterB_n_30));
DFF_X1 \InputRegisterB_dataOut_reg[5]  (.Q (\registerOutB[5] ), .CK (CTS_n617), .D (InputRegisterB_n_29));
DFF_X1 \InputRegisterB_dataOut_reg[6]  (.Q (\registerOutB[6] ), .CK (CTS_n617), .D (InputRegisterB_n_28));
DFF_X1 \InputRegisterB_dataOut_reg[7]  (.Q (\registerOutB[7] ), .CK (CTS_n617), .D (InputRegisterB_n_27));
DFF_X1 \InputRegisterB_dataOut_reg[8]  (.Q (\registerOutB[8] ), .CK (CTS_n617), .D (InputRegisterB_n_26));
DFF_X1 \InputRegisterB_dataOut_reg[9]  (.Q (\registerOutB[9] ), .CK (CTS_n617), .D (InputRegisterB_n_25));
DFF_X1 \InputRegisterB_dataOut_reg[10]  (.Q (\registerOutB[10] ), .CK (CTS_n618), .D (InputRegisterB_n_24));
DFF_X1 \InputRegisterB_dataOut_reg[11]  (.Q (\registerOutB[11] ), .CK (CTS_n618), .D (InputRegisterB_n_23));
DFF_X1 \InputRegisterB_dataOut_reg[12]  (.Q (\registerOutB[12] ), .CK (CTS_n617), .D (InputRegisterB_n_22));
DFF_X1 \InputRegisterB_dataOut_reg[13]  (.Q (\registerOutB[13] ), .CK (CTS_n617), .D (InputRegisterB_n_21));
DFF_X1 \InputRegisterB_dataOut_reg[14]  (.Q (\registerOutB[14] ), .CK (CTS_n618), .D (InputRegisterB_n_20));
DFF_X1 \InputRegisterB_dataOut_reg[15]  (.Q (\registerOutB[15] ), .CK (CTS_n618), .D (InputRegisterB_n_19));
DFF_X1 \InputRegisterB_dataOut_reg[16]  (.Q (\registerOutB[16] ), .CK (CTS_n618), .D (InputRegisterB_n_18));
DFF_X1 \InputRegisterB_dataOut_reg[17]  (.Q (\registerOutB[17] ), .CK (CTS_n618), .D (InputRegisterB_n_17));
DFF_X1 \InputRegisterB_dataOut_reg[18]  (.Q (\registerOutB[18] ), .CK (CTS_n619), .D (InputRegisterB_n_16));
DFF_X1 \InputRegisterB_dataOut_reg[19]  (.Q (\registerOutB[19] ), .CK (CTS_n618), .D (InputRegisterB_n_15));
DFF_X1 \InputRegisterB_dataOut_reg[20]  (.Q (\registerOutB[20] ), .CK (CTS_n619), .D (InputRegisterB_n_14));
DFF_X1 \InputRegisterB_dataOut_reg[21]  (.Q (\registerOutB[21] ), .CK (CTS_n619), .D (InputRegisterB_n_13));
DFF_X1 \InputRegisterB_dataOut_reg[22]  (.Q (\registerOutB[22] ), .CK (CTS_n618), .D (InputRegisterB_n_12));
DFF_X1 \InputRegisterB_dataOut_reg[23]  (.Q (\registerOutB[23] ), .CK (CTS_n619), .D (InputRegisterB_n_11));
DFF_X1 \InputRegisterB_dataOut_reg[24]  (.Q (\registerOutB[24] ), .CK (CTS_n618), .D (InputRegisterB_n_10));
DFF_X1 \InputRegisterB_dataOut_reg[25]  (.Q (\registerOutB[25] ), .CK (CTS_n618), .D (InputRegisterB_n_9));
DFF_X1 \InputRegisterB_dataOut_reg[26]  (.Q (\registerOutB[26] ), .CK (CTS_n618), .D (InputRegisterB_n_8));
DFF_X1 \InputRegisterB_dataOut_reg[27]  (.Q (\registerOutB[27] ), .CK (CTS_n619), .D (InputRegisterB_n_7));
DFF_X1 \InputRegisterB_dataOut_reg[28]  (.Q (\registerOutB[28] ), .CK (CTS_n619), .D (InputRegisterB_n_6));
DFF_X1 \InputRegisterB_dataOut_reg[29]  (.Q (\registerOutB[29] ), .CK (CTS_n617), .D (InputRegisterB_n_5));
DFF_X1 \InputRegisterB_dataOut_reg[30]  (.Q (\registerOutB[30] ), .CK (CTS_n617), .D (InputRegisterB_n_4));
DFF_X1 \InputRegisterB_dataOut_reg[31]  (.Q (\registerOutB[31] ), .CK (CTS_n619), .D (InputRegisterB_n_2));
DFFR_X1 \InputRegisterB_register_reg[0]  (.Q (\InputRegisterB_register[0] ), .CK (CTS_n560)
    , .D (Multiplier[0]), .RN (InputRegisterB_n_1));
DFFR_X1 \InputRegisterB_register_reg[1]  (.Q (\InputRegisterB_register[1] ), .CK (CTS_n560)
    , .D (Multiplier[1]), .RN (InputRegisterB_n_1));
DFFR_X1 \InputRegisterB_register_reg[2]  (.Q (\InputRegisterB_register[2] ), .CK (CTS_n560)
    , .D (Multiplier[2]), .RN (InputRegisterB_n_1));
DFFR_X1 \InputRegisterB_register_reg[3]  (.Q (\InputRegisterB_register[3] ), .CK (CTS_n560)
    , .D (Multiplier[3]), .RN (InputRegisterB_n_1));
DFFR_X1 \InputRegisterB_register_reg[4]  (.Q (\InputRegisterB_register[4] ), .CK (CTS_n560)
    , .D (Multiplier[4]), .RN (InputRegisterB_n_1));
DFFR_X1 \InputRegisterB_register_reg[5]  (.Q (\InputRegisterB_register[5] ), .CK (CTS_n560)
    , .D (Multiplier[5]), .RN (InputRegisterB_n_1));
DFFR_X1 \InputRegisterB_register_reg[6]  (.Q (\InputRegisterB_register[6] ), .CK (CTS_n560)
    , .D (Multiplier[6]), .RN (InputRegisterB_n_1));
DFFR_X1 \InputRegisterB_register_reg[7]  (.Q (\InputRegisterB_register[7] ), .CK (CTS_n560)
    , .D (Multiplier[7]), .RN (InputRegisterB_n_1));
DFFR_X1 \InputRegisterB_register_reg[8]  (.Q (\InputRegisterB_register[8] ), .CK (CTS_n560)
    , .D (Multiplier[8]), .RN (InputRegisterB_n_1));
DFFR_X1 \InputRegisterB_register_reg[9]  (.Q (\InputRegisterB_register[9] ), .CK (CTS_n560)
    , .D (Multiplier[9]), .RN (InputRegisterB_n_1));
DFFR_X1 \InputRegisterB_register_reg[10]  (.Q (\InputRegisterB_register[10] ), .CK (CTS_n560)
    , .D (Multiplier[10]), .RN (InputRegisterB_n_1));
DFFR_X1 \InputRegisterB_register_reg[11]  (.Q (\InputRegisterB_register[11] ), .CK (CTS_n560)
    , .D (Multiplier[11]), .RN (InputRegisterB_n_1));
DFFR_X1 \InputRegisterB_register_reg[12]  (.Q (\InputRegisterB_register[12] ), .CK (CTS_n560)
    , .D (Multiplier[12]), .RN (InputRegisterB_n_1));
DFFR_X1 \InputRegisterB_register_reg[13]  (.Q (\InputRegisterB_register[13] ), .CK (CTS_n560)
    , .D (Multiplier[13]), .RN (InputRegisterB_n_1));
DFFR_X1 \InputRegisterB_register_reg[14]  (.Q (\InputRegisterB_register[14] ), .CK (CTS_n560)
    , .D (Multiplier[14]), .RN (InputRegisterB_n_1));
DFFR_X1 \InputRegisterB_register_reg[15]  (.Q (\InputRegisterB_register[15] ), .CK (CTS_n560)
    , .D (Multiplier[15]), .RN (InputRegisterB_n_1));
DFFR_X1 \InputRegisterB_register_reg[16]  (.Q (\InputRegisterB_register[16] ), .CK (CTS_n560)
    , .D (Multiplier[16]), .RN (InputRegisterB_n_1));
DFFR_X1 \InputRegisterB_register_reg[17]  (.Q (\InputRegisterB_register[17] ), .CK (CTS_n560)
    , .D (Multiplier[17]), .RN (InputRegisterB_n_1));
DFFR_X1 \InputRegisterB_register_reg[18]  (.Q (\InputRegisterB_register[18] ), .CK (CTS_n560)
    , .D (Multiplier[18]), .RN (InputRegisterB_n_1));
DFFR_X1 \InputRegisterB_register_reg[19]  (.Q (\InputRegisterB_register[19] ), .CK (CTS_n560)
    , .D (Multiplier[19]), .RN (InputRegisterB_n_1));
DFFR_X1 \InputRegisterB_register_reg[20]  (.Q (\InputRegisterB_register[20] ), .CK (CTS_n560)
    , .D (Multiplier[20]), .RN (InputRegisterB_n_1));
DFFR_X1 \InputRegisterB_register_reg[21]  (.Q (\InputRegisterB_register[21] ), .CK (CTS_n560)
    , .D (Multiplier[21]), .RN (InputRegisterB_n_1));
DFFR_X1 \InputRegisterB_register_reg[22]  (.Q (\InputRegisterB_register[22] ), .CK (CTS_n560)
    , .D (Multiplier[22]), .RN (InputRegisterB_n_1));
DFFR_X1 \InputRegisterB_register_reg[23]  (.Q (\InputRegisterB_register[23] ), .CK (CTS_n560)
    , .D (Multiplier[23]), .RN (InputRegisterB_n_1));
DFFR_X1 \InputRegisterB_register_reg[24]  (.Q (\InputRegisterB_register[24] ), .CK (CTS_n560)
    , .D (Multiplier[24]), .RN (InputRegisterB_n_1));
DFFR_X1 \InputRegisterB_register_reg[25]  (.Q (\InputRegisterB_register[25] ), .CK (CTS_n560)
    , .D (Multiplier[25]), .RN (InputRegisterB_n_1));
DFFR_X1 \InputRegisterB_register_reg[26]  (.Q (\InputRegisterB_register[26] ), .CK (CTS_n560)
    , .D (Multiplier[26]), .RN (InputRegisterB_n_1));
DFFR_X1 \InputRegisterB_register_reg[27]  (.Q (\InputRegisterB_register[27] ), .CK (CTS_n560)
    , .D (Multiplier[27]), .RN (InputRegisterB_n_1));
DFFR_X1 \InputRegisterB_register_reg[28]  (.Q (\InputRegisterB_register[28] ), .CK (CTS_n560)
    , .D (Multiplier[28]), .RN (InputRegisterB_n_1));
DFFR_X1 \InputRegisterB_register_reg[29]  (.Q (\InputRegisterB_register[29] ), .CK (CTS_n560)
    , .D (Multiplier[29]), .RN (InputRegisterB_n_1));
DFFR_X1 \InputRegisterB_register_reg[30]  (.Q (\InputRegisterB_register[30] ), .CK (CTS_n560)
    , .D (Multiplier[30]), .RN (InputRegisterB_n_1));
DFFR_X1 \InputRegisterB_register_reg[31]  (.Q (\InputRegisterB_register[31] ), .CK (CTS_n560)
    , .D (Multiplier[31]), .RN (InputRegisterB_n_1));
CLKGATETST_X8 InputRegisterB_clk_gate_register_reg (.GCK (CTS_n560), .CK (CTS_n633)
    , .E (enableB), .SE (VSS));
DFF_X1 \InputRegisterA_dataOut_reg[0]  (.Q (slo__n236), .CK (CTS_n618), .D (InputRegisterA_n_34));
DFF_X1 \InputRegisterA_dataOut_reg[1]  (.Q (slo__n198), .CK (CTS_n618), .D (InputRegisterA_n_33));
DFF_X1 \InputRegisterA_dataOut_reg[2]  (.Q (\registerOutA[2] ), .CK (CTS_n618), .D (InputRegisterA_n_32));
DFF_X1 \InputRegisterA_dataOut_reg[3]  (.Q (\registerOutA[3] ), .CK (CTS_n618), .D (InputRegisterA_n_31));
DFF_X1 \InputRegisterA_dataOut_reg[4]  (.Q (\registerOutA[4] ), .CK (CTS_n618), .D (InputRegisterA_n_30));
DFF_X1 \InputRegisterA_dataOut_reg[5]  (.Q (\registerOutA[5] ), .CK (CTS_n618), .D (InputRegisterA_n_29));
DFF_X1 \InputRegisterA_dataOut_reg[6]  (.Q (\registerOutA[6] ), .CK (CTS_n618), .D (InputRegisterA_n_28));
DFF_X1 \InputRegisterA_dataOut_reg[7]  (.Q (\registerOutA[7] ), .CK (CTS_n618), .D (InputRegisterA_n_27));
DFF_X1 \InputRegisterA_dataOut_reg[8]  (.Q (\registerOutA[8] ), .CK (CTS_n617), .D (InputRegisterA_n_26));
DFF_X1 \InputRegisterA_dataOut_reg[9]  (.Q (\registerOutA[9] ), .CK (CTS_n617), .D (InputRegisterA_n_25));
DFF_X1 \InputRegisterA_dataOut_reg[10]  (.Q (\registerOutA[10] ), .CK (CTS_n617), .D (InputRegisterA_n_24));
DFF_X1 \InputRegisterA_dataOut_reg[11]  (.Q (\registerOutA[11] ), .CK (CTS_n617), .D (InputRegisterA_n_23));
DFF_X1 \InputRegisterA_dataOut_reg[12]  (.Q (\registerOutA[12] ), .CK (CTS_n617), .D (InputRegisterA_n_22));
DFF_X1 \InputRegisterA_dataOut_reg[13]  (.Q (\registerOutA[13] ), .CK (CTS_n617), .D (InputRegisterA_n_21));
DFF_X1 \InputRegisterA_dataOut_reg[14]  (.Q (\registerOutA[14] ), .CK (CTS_n617), .D (InputRegisterA_n_20));
DFF_X1 \InputRegisterA_dataOut_reg[15]  (.Q (\registerOutA[15] ), .CK (CTS_n617), .D (InputRegisterA_n_19));
DFF_X1 \InputRegisterA_dataOut_reg[16]  (.Q (\registerOutA[16] ), .CK (CTS_n617), .D (InputRegisterA_n_18));
DFF_X1 \InputRegisterA_dataOut_reg[17]  (.Q (\registerOutA[17] ), .CK (CTS_n617), .D (InputRegisterA_n_17));
DFF_X1 \InputRegisterA_dataOut_reg[18]  (.Q (\registerOutA[18] ), .CK (CTS_n617), .D (InputRegisterA_n_16));
DFF_X1 \InputRegisterA_dataOut_reg[19]  (.Q (\registerOutA[19] ), .CK (CTS_n617), .D (InputRegisterA_n_15));
DFF_X1 \InputRegisterA_dataOut_reg[20]  (.Q (\registerOutA[20] ), .CK (CTS_n617), .D (InputRegisterA_n_14));
DFF_X1 \InputRegisterA_dataOut_reg[21]  (.Q (\registerOutA[21] ), .CK (CTS_n617), .D (InputRegisterA_n_13));
DFF_X1 \InputRegisterA_dataOut_reg[22]  (.Q (\registerOutA[22] ), .CK (CTS_n617), .D (InputRegisterA_n_12));
DFF_X1 \InputRegisterA_dataOut_reg[23]  (.Q (\registerOutA[23] ), .CK (CTS_n619), .D (InputRegisterA_n_11));
DFF_X1 \InputRegisterA_dataOut_reg[24]  (.Q (\registerOutA[24] ), .CK (CTS_n617), .D (InputRegisterA_n_10));
DFF_X1 \InputRegisterA_dataOut_reg[25]  (.Q (\registerOutA[25] ), .CK (CTS_n619), .D (InputRegisterA_n_9));
DFF_X1 \InputRegisterA_dataOut_reg[26]  (.Q (\registerOutA[26] ), .CK (CTS_n619), .D (InputRegisterA_n_8));
DFF_X1 \InputRegisterA_dataOut_reg[27]  (.Q (\registerOutA[27] ), .CK (CTS_n619), .D (InputRegisterA_n_7));
DFF_X1 \InputRegisterA_dataOut_reg[28]  (.Q (\registerOutA[28] ), .CK (CTS_n618), .D (InputRegisterA_n_6));
DFF_X1 \InputRegisterA_dataOut_reg[29]  (.Q (\registerOutA[29] ), .CK (CTS_n618), .D (InputRegisterA_n_5));
DFF_X1 \InputRegisterA_dataOut_reg[30]  (.Q (\registerOutA[30] ), .CK (CTS_n619), .D (InputRegisterA_n_4));
DFF_X1 \InputRegisterA_dataOut_reg[31]  (.Q (\registerOutA[31] ), .CK (CTS_n618), .D (InputRegisterA_n_2));
DFFR_X1 \InputRegisterA_register_reg[0]  (.Q (\InputRegisterA_register[0] ), .CK (CTS_n564)
    , .D (CLOCK_slh_n870), .RN (InputRegisterA_n_1));
DFFR_X1 \InputRegisterA_register_reg[1]  (.Q (\InputRegisterA_register[1] ), .CK (CTS_n564)
    , .D (CLOCK_slh_n840), .RN (InputRegisterA_n_1));
DFFR_X1 \InputRegisterA_register_reg[2]  (.Q (\InputRegisterA_register[2] ), .CK (CTS_n564)
    , .D (Multiplicand[2]), .RN (InputRegisterA_n_1));
DFFR_X1 \InputRegisterA_register_reg[3]  (.Q (\InputRegisterA_register[3] ), .CK (CTS_n564)
    , .D (sph_n1162), .RN (InputRegisterA_n_1));
DFFR_X1 \InputRegisterA_register_reg[4]  (.Q (\InputRegisterA_register[4] ), .CK (CTS_n564)
    , .D (sph__n1163), .RN (InputRegisterA_n_1));
DFFR_X1 \InputRegisterA_register_reg[5]  (.Q (\InputRegisterA_register[5] ), .CK (CTS_n564)
    , .D (Multiplicand[5]), .RN (InputRegisterA_n_1));
DFFR_X1 \InputRegisterA_register_reg[6]  (.Q (\InputRegisterA_register[6] ), .CK (CTS_n564)
    , .D (Multiplicand[6]), .RN (InputRegisterA_n_1));
DFFR_X1 \InputRegisterA_register_reg[7]  (.Q (\InputRegisterA_register[7] ), .CK (CTS_n564)
    , .D (sph_n1154), .RN (InputRegisterA_n_1));
DFFR_X1 \InputRegisterA_register_reg[8]  (.Q (\InputRegisterA_register[8] ), .CK (CTS_n564)
    , .D (sph_n1217), .RN (InputRegisterA_n_1));
DFFR_X1 \InputRegisterA_register_reg[9]  (.Q (\InputRegisterA_register[9] ), .CK (CTS_n564)
    , .D (sph__n1207), .RN (InputRegisterA_n_1));
DFFR_X1 \InputRegisterA_register_reg[10]  (.Q (\InputRegisterA_register[10] ), .CK (CTS_n564)
    , .D (sph__n1195), .RN (InputRegisterA_n_1));
DFFR_X1 \InputRegisterA_register_reg[11]  (.Q (\InputRegisterA_register[11] ), .CK (CTS_n564)
    , .D (CLOCK_slh_n928), .RN (InputRegisterA_n_1));
DFFR_X1 \InputRegisterA_register_reg[12]  (.Q (\InputRegisterA_register[12] ), .CK (CTS_n564)
    , .D (sph__n1201), .RN (InputRegisterA_n_1));
DFFR_X1 \InputRegisterA_register_reg[13]  (.Q (\InputRegisterA_register[13] ), .CK (CTS_n564)
    , .D (sph_n1182), .RN (InputRegisterA_n_1));
DFFR_X1 \InputRegisterA_register_reg[14]  (.Q (\InputRegisterA_register[14] ), .CK (CTS_n564)
    , .D (sph__n1192), .RN (InputRegisterA_n_1));
DFFR_X1 \InputRegisterA_register_reg[15]  (.Q (\InputRegisterA_register[15] ), .CK (CTS_n564)
    , .D (sph__n1198), .RN (InputRegisterA_n_1));
DFFR_X1 \InputRegisterA_register_reg[16]  (.Q (\InputRegisterA_register[16] ), .CK (CTS_n564)
    , .D (sph__n1169), .RN (InputRegisterA_n_1));
DFFR_X1 \InputRegisterA_register_reg[17]  (.Q (\InputRegisterA_register[17] ), .CK (CTS_n564)
    , .D (sph__n1166), .RN (InputRegisterA_n_1));
DFFR_X1 \InputRegisterA_register_reg[18]  (.Q (\InputRegisterA_register[18] ), .CK (CTS_n564)
    , .D (sph__n1204), .RN (InputRegisterA_n_1));
DFFR_X1 \InputRegisterA_register_reg[19]  (.Q (\InputRegisterA_register[19] ), .CK (CTS_n564)
    , .D (CLOCK_slh__n943), .RN (InputRegisterA_n_1));
DFFR_X1 \InputRegisterA_register_reg[20]  (.Q (\InputRegisterA_register[20] ), .CK (CTS_n564)
    , .D (sph__n1189), .RN (InputRegisterA_n_1));
DFFR_X1 \InputRegisterA_register_reg[21]  (.Q (\InputRegisterA_register[21] ), .CK (CTS_n564)
    , .D (sph__n1186), .RN (InputRegisterA_n_1));
DFFR_X1 \InputRegisterA_register_reg[22]  (.Q (\InputRegisterA_register[22] ), .CK (CTS_n564)
    , .D (sph__n1172), .RN (InputRegisterA_n_1));
DFFR_X1 \InputRegisterA_register_reg[23]  (.Q (\InputRegisterA_register[23] ), .CK (CTS_n565)
    , .D (Multiplicand[23]), .RN (InputRegisterA_n_1));
DFFR_X1 \InputRegisterA_register_reg[24]  (.Q (\InputRegisterA_register[24] ), .CK (CTS_n564)
    , .D (sph__n1183), .RN (InputRegisterA_n_1));
DFFR_X1 \InputRegisterA_register_reg[25]  (.Q (\InputRegisterA_register[25] ), .CK (CTS_n565)
    , .D (sph__n1144), .RN (InputRegisterA_n_1));
DFFR_X1 \InputRegisterA_register_reg[26]  (.Q (\InputRegisterA_register[26] ), .CK (CTS_n565)
    , .D (sph__n1141), .RN (InputRegisterA_n_1));
DFFR_X1 \InputRegisterA_register_reg[27]  (.Q (\InputRegisterA_register[27] ), .CK (CTS_n565)
    , .D (Multiplicand[27]), .RN (InputRegisterA_n_1));
DFFR_X1 \InputRegisterA_register_reg[28]  (.Q (\InputRegisterA_register[28] ), .CK (CTS_n564)
    , .D (CLOCK_slh_n845), .RN (InputRegisterA_n_1));
DFFR_X1 \InputRegisterA_register_reg[29]  (.Q (\InputRegisterA_register[29] ), .CK (CTS_n565)
    , .D (CLOCK_slh_n800), .RN (InputRegisterA_n_1));
DFFR_X1 \InputRegisterA_register_reg[30]  (.Q (\InputRegisterA_register[30] ), .CK (CTS_n565)
    , .D (sph_n1140), .RN (InputRegisterA_n_1));
DFFR_X1 \InputRegisterA_register_reg[31]  (.Q (\InputRegisterA_register[31] ), .CK (CTS_n565)
    , .D (CLOCK_slh_n790), .RN (InputRegisterA_n_1));
CLKGATETST_X8 InputRegisterA_clk_gate_register_reg (.GCK (CTS_n602), .CK (CTS_n633)
    , .E (hfn_ipo_n72), .SE (VSS));
BoothAlgorithmMultiplier BAMMultiplier (.Product ({\registerInProduct[63] , \registerInProduct[62] , 
    \registerInProduct[61] , \registerInProduct[60] , \registerInProduct[59] , \registerInProduct[58] , 
    \registerInProduct[57] , \registerInProduct[56] , \registerInProduct[55] , \registerInProduct[54] , 
    \registerInProduct[53] , \registerInProduct[52] , \registerInProduct[51] , \registerInProduct[50] , 
    \registerInProduct[49] , \registerInProduct[48] , \registerInProduct[47] , \registerInProduct[46] , 
    \registerInProduct[45] , \registerInProduct[44] , \registerInProduct[43] , \registerInProduct[42] , 
    \registerInProduct[41] , \registerInProduct[40] , \registerInProduct[39] , \registerInProduct[38] , 
    \registerInProduct[37] , \registerInProduct[36] , \registerInProduct[35] , \registerInProduct[34] , 
    \registerInProduct[33] , \registerInProduct[32] , \registerInProduct[31] , \registerInProduct[30] , 
    \registerInProduct[29] , \registerInProduct[28] , \registerInProduct[27] , \registerInProduct[26] , 
    \registerInProduct[25] , \registerInProduct[24] , \registerInProduct[23] , \registerInProduct[22] , 
    \registerInProduct[21] , \registerInProduct[20] , \registerInProduct[19] , \registerInProduct[18] , 
    \registerInProduct[17] , \registerInProduct[16] , \registerInProduct[15] , \registerInProduct[14] , 
    \registerInProduct[13] , \registerInProduct[12] , \registerInProduct[11] , \registerInProduct[10] , 
    \registerInProduct[9] , \registerInProduct[8] , \registerInProduct[7] , \registerInProduct[6] , 
    \registerInProduct[5] , \registerInProduct[4] , \registerInProduct[3] , \registerInProduct[2] , 
    \registerInProduct[1] , \registerInProduct[0] }), .Multiplicand ({\registerOutA[31] , 
    \registerOutA[30] , \registerOutA[29] , \registerOutA[28] , \registerOutA[27] , 
    \registerOutA[26] , \registerOutA[25] , \registerOutA[24] , \registerOutA[23] , 
    \registerOutA[22] , \registerOutA[21] , \registerOutA[20] , \registerOutA[19] , 
    \registerOutA[18] , \registerOutA[17] , \registerOutA[16] , \registerOutA[15] , 
    \registerOutA[14] , \registerOutA[13] , \registerOutA[12] , \registerOutA[11] , 
    \registerOutA[10] , \registerOutA[9] , \registerOutA[8] , \registerOutA[7] , 
    \registerOutA[6] , \registerOutA[5] , \registerOutA[4] , \registerOutA[3] , \registerOutA[2] , 
    slo__n198, slo__n236}), .Multiplier ({drc_ipo_n105, \registerOutB[30] , drc_ipo_n104, 
    drc_ipo_n103, drc_ipo_n102, drc_ipo_n354, drc_ipo_n100, drc_ipo_n99, drc_ipo_n98, 
    drc_ipo_n97, drc_ipo_n96, drc_ipo_n95, drc_ipo_n94, drc_ipo_n93, drc_ipo_n92, 
    drc_ipo_n91, drc_ipo_n90, drc_ipo_n89, drc_ipo_n88, drc_ipo_n87, drc_ipo_n86, 
    drc_ipo_n85, drc_ipo_n84, drc_ipo_n83, drc_ipo_n82, \registerOutB[6] , drc_ipo_n80, 
    drc_ipo_n79, drc_ipo_n78, \registerOutB[2] , drc_ipo_n76, opt_ipo_n299}), .Multiplier_0_PP_0 (opt_ipo_n299)
    , .drc_ipoPP_0 (drc_ipo_n347), .drc_ipoPP_1 (drc_ipo_n348), .drc_ipoPP_2 (drc_ipo_n88)
    , .drc_ipoPP_3 (drc_ipo_n350), .drc_ipoPP_4 (drc_ipo_n351), .drc_ipoPP_5 (drc_ipo_n352)
    , .drc_ipoPP_6 (drc_ipo_n353), .drc_ipoPP_7 (drc_ipo_n355), .Multiplier_19_PP_2 (drc_ipo_n94)
    , .drc_ipoPP_3PP_0 (drc_ipo_n350), .drc_ipoPP_2PP_0 (drc_ipo_n88));
BUF_X32 hfn_ipo_c71 (.Z (hfn_ipo_n71), .A (enableA));
BUF_X2 hfn_ipo_c72 (.Z (hfn_ipo_n72), .A (enableA));
BUF_X32 drc_ipo_c356 (.Z (drc_ipo_n347), .A (drc_ipo_n83));
BUF_X8 hfn_ipo_c74 (.Z (hfn_ipo_n74), .A (OutputRegister_n_1));
BUF_X16 drc_ipo_c105 (.Z (drc_ipo_n105), .A (\registerOutB[31] ));
BUF_X16 drc_ipo_c104 (.Z (drc_ipo_n104), .A (\registerOutB[29] ));
BUF_X32 drc_ipo_c103 (.Z (drc_ipo_n103), .A (\registerOutB[28] ));
BUF_X32 drc_ipo_c102 (.Z (drc_ipo_n102), .A (\registerOutB[27] ));
BUF_X32 drc_ipo_c101 (.Z (drc_ipo_n101), .A (\registerOutB[26] ));
BUF_X32 drc_ipo_c100 (.Z (drc_ipo_n100), .A (\registerOutB[25] ));
BUF_X32 drc_ipo_c99 (.Z (drc_ipo_n99), .A (\registerOutB[24] ));
BUF_X32 drc_ipo_c98 (.Z (drc_ipo_n98), .A (\registerOutB[23] ));
BUF_X32 drc_ipo_c97 (.Z (drc_ipo_n97), .A (\registerOutB[22] ));
BUF_X32 drc_ipo_c96 (.Z (drc_ipo_n96), .A (\registerOutB[21] ));
BUF_X32 drc_ipo_c95 (.Z (drc_ipo_n95), .A (\registerOutB[20] ));
BUF_X16 drc_ipo_c94 (.Z (drc_ipo_n94), .A (\registerOutB[19] ));
BUF_X32 drc_ipo_c93 (.Z (drc_ipo_n93), .A (\registerOutB[18] ));
BUF_X32 drc_ipo_c92 (.Z (drc_ipo_n92), .A (\registerOutB[17] ));
BUF_X8 drc_ipo_c91 (.Z (drc_ipo_n91), .A (\registerOutB[16] ));
BUF_X16 drc_ipo_c90 (.Z (drc_ipo_n90), .A (\registerOutB[15] ));
BUF_X32 drc_ipo_c89 (.Z (drc_ipo_n89), .A (\registerOutB[14] ));
BUF_X8 drc_ipo_c88 (.Z (drc_ipo_n88), .A (\registerOutB[13] ));
BUF_X16 drc_ipo_c87 (.Z (drc_ipo_n87), .A (\registerOutB[12] ));
BUF_X32 drc_ipo_c86 (.Z (drc_ipo_n86), .A (\registerOutB[11] ));
BUF_X32 drc_ipo_c85 (.Z (drc_ipo_n85), .A (\registerOutB[10] ));
BUF_X32 drc_ipo_c84 (.Z (drc_ipo_n84), .A (\registerOutB[9] ));
BUF_X32 drc_ipo_c83 (.Z (drc_ipo_n83), .A (\registerOutB[8] ));
BUF_X16 drc_ipo_c82 (.Z (drc_ipo_n82), .A (\registerOutB[7] ));
CLKBUF_X1 CLOCK_slh__c755 (.Z (CLOCK_slh_n790), .A (Multiplicand[31]));
BUF_X2 drc_ipo_c80 (.Z (drc_ipo_n80), .A (\registerOutB[5] ));
BUF_X16 drc_ipo_c79 (.Z (drc_ipo_n79), .A (\registerOutB[4] ));
BUF_X16 drc_ipo_c78 (.Z (drc_ipo_n78), .A (\registerOutB[3] ));
BUF_X32 drc_ipo_c360 (.Z (drc_ipo_n351), .A (drc_ipo_n92));
BUF_X4 drc_ipo_c76 (.Z (drc_ipo_n76), .A (\registerOutB[1] ));
BUF_X32 drc_ipo_c362 (.Z (drc_ipo_n353), .A (drc_ipo_n101));
BUF_X4 drc_ipo_c363 (.Z (drc_ipo_n354), .A (drc_ipo_n101));
INV_X8 CTS_L6_c575 (.ZN (CTS_n565), .A (CTS_n603));
CLKBUF_X1 sph__c1029 (.Z (sph_n1140), .A (Multiplicand[30]));
BUF_X8 opt_ipo_c308 (.Z (opt_ipo_n299), .A (slo___n231));
BUF_X32 drc_ipo_c361 (.Z (drc_ipo_n352), .A (drc_ipo_n98));
INV_X8 CTS_L6_c611 (.ZN (CTS_n619), .A (CTS_n630));
BUF_X32 drc_ipo_c357 (.Z (drc_ipo_n348), .A (drc_ipo_n84));
BUF_X8 drc_ipo_c359 (.Z (drc_ipo_n350), .A (drc_ipo_n91));
BUF_X32 drc_ipo_c364 (.Z (drc_ipo_n355), .A (drc_ipo_n102));
INV_X32 CTS_L4_c625 (.ZN (CTS_n631), .A (CTS_n633));
BUF_X8 CTS_L1_c671 (.Z (CTS_n707), .A (clk));
INV_X8 CTS_L5_c622 (.ZN (CTS_n630), .A (CTS_n631));
INV_X8 CTS_L6_c574 (.ZN (CTS_n564), .A (CTS_n603));
CLKBUF_X1 CLOCK_slh__c759 (.Z (CLOCK_slh_n800), .A (Multiplicand[29]));
INV_X16 CTS_L6_c610 (.ZN (CTS_n618), .A (CTS_n630));
INV_X8 CTS_L5_c602 (.ZN (CTS_n603), .A (CTS_n602));
INV_X8 CTS_L3_c632 (.ZN (CTS_n633), .A (CTS_n634));
INV_X4 CTS_L2_c635 (.ZN (CTS_n634), .A (CTS_n707));
CLKBUF_X1 sph__c1032 (.Z (sph__n1141), .A (Multiplicand[26]));
CLKBUF_X1 sph__c1035 (.Z (sph__n1144), .A (Multiplicand[25]));
CLKBUF_X1 sph__c1038 (.Z (sph_n1154), .A (Multiplicand[7]));
CLKBUF_X1 sph__c1041 (.Z (sph_n1162), .A (Multiplicand[3]));
CLKBUF_X1 sph__c1044 (.Z (sph__n1163), .A (Multiplicand[4]));
CLKBUF_X1 sph__c1047 (.Z (sph__n1166), .A (Multiplicand[17]));
CLKBUF_X1 sph__c1050 (.Z (sph__n1169), .A (Multiplicand[16]));
CLKBUF_X1 CLOCK_slh__c775 (.Z (CLOCK_slh_n840), .A (Multiplicand[1]));
CLKBUF_X1 CLOCK_slh__c777 (.Z (CLOCK_slh_n845), .A (Multiplicand[28]));
CLKBUF_X1 sph__c1053 (.Z (sph__n1172), .A (Multiplicand[22]));
CLKBUF_X1 sph__c1056 (.Z (sph_n1182), .A (Multiplicand[13]));
CLKBUF_X1 sph__c1059 (.Z (sph__n1183), .A (Multiplicand[24]));
CLKBUF_X1 sph__c1062 (.Z (sph__n1186), .A (Multiplicand[21]));
CLKBUF_X1 CLOCK_slh__c787 (.Z (CLOCK_slh_n870), .A (Multiplicand[0]));
CLKBUF_X1 sph__c1065 (.Z (sph__n1189), .A (Multiplicand[20]));
CLKBUF_X1 sph__c1068 (.Z (sph__n1192), .A (Multiplicand[14]));
CLKBUF_X1 sph__c1071 (.Z (sph__n1195), .A (Multiplicand[10]));
CLKBUF_X1 sph__c1074 (.Z (sph__n1198), .A (Multiplicand[15]));
CLKBUF_X1 sph__c1077 (.Z (sph__n1201), .A (Multiplicand[12]));
CLKBUF_X1 sph__c1080 (.Z (sph__n1204), .A (Multiplicand[18]));
CLKBUF_X1 sph__c1083 (.Z (sph__n1207), .A (Multiplicand[9]));
CLKBUF_X1 sph__c1086 (.Z (sph_n1217), .A (Multiplicand[8]));
CLKBUF_X1 CLOCK_slh__c812 (.Z (CLOCK_slh_n928), .A (Multiplicand[11]));
CLKBUF_X1 CLOCK_slh__c820 (.Z (CLOCK_slh__n943), .A (Multiplicand[19]));
CLKBUF_X2 CLOCK_spc__L1_c894 (.Z (CLOCK_spc__n1018), .A (OutputRegister_n_1));

endmodule //BAMIntegrated


