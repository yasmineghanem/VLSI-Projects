module SequentialMultiplier ();
    
endmodule